BZh91AY&SY�B�A 	_�Py���g߰����`�8��  �t
TP����i�  h    �=�cJJ��ѧ��	��bh� ���U44M���  5=4"� � 4d   ���a2dɑ��4�# C �!!�d�I��ѽS  ��M3�H>�$���^# �����D�Џ�@(���f��B�E,�,n�&Kb���n�=��ȭ�$
 ( AP@��L�ҵ���( �+"��QI4��D!쐌�R�K�K���"�q^B%�c]ŋ���2��Ln=��f�(M!�;U�<	VD�A��C=�9�Ob�\�v�#�<����n҆�Q�_t�����h��� A+��&,2�ϛ'�I��v:�es`�m���o9m���M��fEݼ̼m�l�ۖ�'33'o���a��n��uխkJֲ����� �c~���j�y�<�G��>A狟C��uk��4�0db�["�y��I&���`�{��W�8��$FW^�ڸ4Z��J�a����p��x�:뮑�8�߁��b	=��!.��9f���\ȑ��R��@�%hd� �F�k��]uF!���*Y$�O�`�C �LD�� x�@�Z�#� \<=�<���b d�fO� �� l�$�I(u:��]	�� hV����&L�Ś�	����6r��mj�� Xњ�7�FQ$�I��p�]��}�pّ���v�+�u�PB�*$u�B�.��K,�:Y�Un���j.fC�(�pp�D��Ww�+�rE��&`;�����r'�7ulHͮ�9d�I&ݙQ,O\�f�t�<��j��m!mR��LQ�	�9�.qH�&�I$�[�3��ȆR�y7���-U^���Q���D<�(ى��8x�I$�J�}�5.�w6mmP��24���Ԍ�Sh��ք.��J#T�RI$���ٶ�u�GD,�Ls\)���?u�v+%(k`O}�`�~P=��{`� 8������%9�Ԥ����"��A �>;�� �� ����l���c0d�c6�L����6��hP�䆼�Hp�r�j�}��BI&Ѐl���H�����9�����;����+x�F�b���g���N���;`���s8���5 ��K^�V.=G���}ʶ���W9���׬S�	@�澥�3�#$�5�>�eB�͔ 0]���0aXz���R�ncA"�3]m��	�2��-����4��ni ��,�FE�x�r>�Z�&�0U]A`S"��l���
�C$ZS�����O��7I z��N�0�o��<��$.zb�9,L��y��|q����䒸� ����x���pݓ�و�cf��ؐ����9>�3M��h*�(�d��s����M! �j� �稁q&���(C�b&+���F�C"ʐAk��9�@B&�V�6�Pv� q�ƨ���T�����onՠ�����`��KI�w�ղŤ D#x�n=]+�� iT=�XP�$fD��Rɐjc�2%�7+-1O�@A���KK�<xJ���� X��3��'GFrM�@���e| i�F�\����*�"�����
��ᩦKE;�K�뉤�f`1(��w$S�	�/�