BZh91AY&SYcԦ$ �_�Px����߰����`�l�  =��̒��	"�����S�Ğ�Oj z�i�6�z ��$�=M�M    �s F	�0M`�L$����F�    Q�A����# �4���0�$�Di1Fi=MO)�6P�= @�i4X��!x)`U$(Y�=o�D��.��O#P<O�	A���!�$N�(-�:#��p�����::h��l���K �28e�Oo_���_�����2@�f	i��C��qÃ�b�-�J��Aj+�=�#������hh�P�'��ʏ^�ԉt�@�P���+L��u��@��<ug�sp�l��3nV,F�`�������AA����<���� |K�4Hi���g�gT��49S��ƾs�A����aE������0�&�[s��^�ٍ{W�5��Z���z�l�em�ڽ����̻���P�)JYK)�#ǧX��#rM�bG�nY�C�d�a�`��v��~�y;���['��Ԉ�D�˫b�Wލ�|���$�WcK8�:�	E.3�0,��$H��^�).}�m�YVe���dtI��H9�1��`�*������-w��
 j�F���z��,h\yN�N0*�\S������*/�����:돠�7�ԋ7��6p<�UԤ��oV���`l>��<}�D���h�����烙]|����zH�o^��* ��U�҅F�7%UkU'�:"��ck�`;@OS@��=�&*�a�߀�s��k���#��:A&�PD��2�����M���6rk#
�]���컾Č�����$�r���%�x{���l�O��[*sb:�'gb����^�,nP7x.-Դ���)J޹*�fY8�sy"�����)���j�Rf�7/"�P{Q�*��U�-(���b��W�uG{}���GeX�o,���ȇ"�{
�9��0���I'�le�I>yl��^z�lEg��frp�<���D�yCu)I.�U�V�T��V�������V��}y�WbDN���"O:2�Т�,om�UW�U���|��+ai ���n���5X���И��C(�A�4(,���DbV���aF�P"`��b*��`��% ~TA������x�VQ"|!��N��0��߸�M�CT5A!B�g��]T�㼨a"Qi����Ѐ�54S�s�7$#٫����o��O�gΛN����Dj�Ν��J���c�P<LC���on�ag�2ĐuH���ǈ�N}�&��m�U�<t��99��?2�<�c�}��'���wof����: �[���.z�bei����}����Pлg�w��u��t6v(���ݍN�h�T@�E'
�Vi�_E��U8��i�fj?��R����V�����@\[�BJ�5�@ߞ/Eq}g͋���HF�\�,������������w��8c��~l2�C�F�9�*�ݏ��lV΂Ff��9p�*�v�+��	"�����O�)�<-!e�t9��Q���-�	� ��c�;)7C����P0�Y1?�R�F���J&�̹���"������V��z�i��(!뤧��j]%ܥ]��-�P[��#��J[�����I����9 ޢ;�%�v��5���ƞ�����Pz�e���J�ک���s�c��Rug�~�:0� Bo�����'Q�ޠ�	@Sk��W���-&\cB�*s5^�a���5�JH�B-q���t�M�w��ԈB�g$P�J-SN���B�"�� !�Q&l����i�4gG����\��_�mj�bB�h"���y�6�+���?���^��UV.�י���H�̎f�+X���3N�:�2:{8�a_���)��1 