BZh91AY&SYSdK ��_�py����߰����`q������*�RD(R���     z  A���U�4��P L@(�vR�顋J� �'�(��� 8�UYb�D�cb Wl�NY$Y���*� �HJ$�ʪ�H�e*���H���Y��J�h ���"�U���B��e$�Yd(�� �*���$U�j@UR	e���+� A �� %*����LL4�a0 "�hĚ��i�     L11�220CFi�F i�# ��H��i�     L10�D�	�4�S�)�x��Ld�OQ��jmF�MA&���F�y �F�  h ���Z���$H�@J��a@E1���$ ��!!�!� ���矤!��ܟ�ɴ�*�'	$� �g���Z�?F� ���C$*!���g��Wl=��g�=�<���P@� ��aE$"�H��XAd X �a�H��d��@@"�$@"���X�(q�H �"� ��$���(B)"�XE 
AHE�(�, )�,���RABE,���
@ RE���)�$��B��(�a �I ��a���o�S�l��_����w���SN��S_�X�7�ov�m�8�ӽ;ѵ�ZG�Zg���)RR�"���r�LA��AU?��U���:E�y�/
2E�P0� �SG S..��R2�Jɢ��eE���@K�I�Xg.I��'1M+���jb�9�p�B�ɹ
�$T����v��9Me����m
m��2rV" ��ə�*�Qx�"��bڨ&�Na����g���J��.��LЛN�ut�d# Ǚ�.�f :��w/��J6p�� �����"�ND�b2��r��wn�4% ���I$��X�A�5���t�d�&�l��C��<�T��̪XY	cI�`ʥ`�Ӄm�A&�c�v���G��Nŵ�L"n(5+21	����M���P�l�q)���-�<�țhT�1�f(�ł�J�D(���D�x
���!eT������^N2&Bu��s��VT����Z�7�����l�S9�\�V�2��b]1QP���B�Y	�S*K��ː�A�J�Z����bm��j����ST�#ffk��Q��C0�2`I�)	T�Ij%d�J�7�ú�7����û�h����!f:��RC ،�%:[�S' �d���!$���-����4lT!f@�9tM # ���R��l���5N@c<���Ab�ZU(�+�	WY���N<���r`6i��$��YF�J��*� ٻ�-�6f���%����O�A�b�d�ك6��a�0	h�*&��M�C�H���-�K�3T�C`)������u+N�t~�S���T���Ȝ��Kg�xg�K��F.*FS
*��U#�OE̅����a٫˚H��/�%���&J�ᠨM�Ż��@0I�4�-���U��M��P?^,�2�\ ���$�y�&EL��y��T���@in��������LI�.�D� e:a�Q5OwS�Ysl�b��.h�a�KH�N�AE�x�P��lUDԅh�7p`Q�)�	�����QG.h j�TD('$A"�`QjY78椪�w.b�&�$"�'Pe��.�b���ab����(�iQ�J�aZ@���؉�*����`�Л�h�-��^tɋ�aၒ��ʓf��C��T]��ؤ͕Urd
�IUc!<�+�os_'N
�"�����f'M&p9��A%
��UD�T���6\ZVҫ�f���kb�C/%d�o);ED̅n�5jr�E�5%	�-�NVL,�X��f�"QZ����(]Rc���	�"f�P,��� ���_6�e6��x�m�uq'�~ ����������8j	����߹����n�b|~Q>������|��%��ef�2��`v��(�ι�l���Ն���K�k)��Ͷ-M)Ivن���1���2L0H�ǈ��A,�a���#�<�]6��1-�+��QXҐ�X��\1�P�]�46���ѭ3nt��:2�d����Xjj�Mu�����ԘI�K���$��Q�����&.�W::�ɍF�)��mJb�]���6-�����[q7�v]���mR�:�SK�^�M�kb�Wg`��t˚�M �q��v��SK*�!.LUP��;�j��h	�s j�\�bR�e LT�M�����rh1v!��#��sF��v�ln͵Sa�kNl1Ոn�#&l�]!3��Z�i5��r�\˰Vf;��q���l��k�r���Hy��xLOθ�UB�k@+PqCe�$6�X5��;;%���dq�Y���3u�r%5��۶��ŕѕ�j8�V�d,D�����&m-��[��l��+�B�5�V���t�l1m!���!r:�AM)h岱
�Q֣0��m�*�,p�\v�:<k^�b�΀E�XZl�Y`�V�f��5Ķ�� f�RZ%0��R�4ua1CF6��]��5��Gm��CLg����iqQ����j����x#v�!�PPVPuѣtU�q���m��F�R�n�^c�njeu��۴[��:�.4�M��WJQ���04�a�ź�$��`ؤ�B�P��e�GZM,��f[l��Yh�D���d��2�kf��Θ&Q�j��X]��8l�5&j��ktM6Bh��LVf��V�k���b�Dg���̗X\Sk��e���m�F`y�+U�u��m�Sb�45ѴQ�W&%�b�V�J�lF�lb\�sĩv��]3�1�ژ�Zݣ�6�K]�e���]u���P��b(��B�:���q�4��F�.�q-IU�n��ku�{K]:̦�5�\���?0BI}!�q��@K,���hL�-Q&��Wb���,�Y	��C�`@YHB�H( ,�B{k$�B)�� �
H)"�U�X)$��IRLH,X���I0�@P�6ɽ�1`��J�Yąd�+&�LHe�Z�$��P�q��|�`T
.o&"ɛ����,d1\CIěC4���6��l5��	�¤ݪ��6͢2f���&��sv;�Xb�S+Gb
,�T16�5VE���,�*�l1�5Ct�N�wt��kX±���Ƥ8�f�9���EA��a*(�M!�XX�x�&��jP4�]:A����q�;�b�,���հY��Ш=�y�^0���"�t�:խ\�E���e�텙eE��Si�M"���5zy�T�l�t��&�4�7l7�ʰU�)�.�SH�.VԻi�4��5�]��Y�^r���LC�S3i]5
�Y��_{����M-�����l���xZt.��S�4�t�t��Zc6��xg9��W()*�x�R�2�S�1:�嗶��B�x\�noNG��76��jT��|f�Q�+��g��d-��7ֳcz���}�����I"
A/3�A�G�:�-���K����zg�l�e'M�t���R�R����(ZVT�~E�U�*��\�06�0m�n,Ma2�acYC���36�
�5u��KBiB�`�0Γc��ҹ�MZ�kiR2[f��%�و��`Vkq,)V.i`�31WI[��c(��C B0BEs���j�[@����SmJ�GEv2Kv�Jd���`�Z8�l�����v�e���K�.bm�kWX�Me�c�e3.��I8�Iɤ|��ƻZ[�!���ȫ�M���e�n�W��$۳CY�i���ba�?���,��d)0:a��t�'{�4����(v�Gn8��J��g_��j�Ci
����|��]+�N�����N٤8�yӀoua�߯�W�*AN�[�`n��|<<뜓X=-�����%`��w�w�Q�2á��2q��h���r�^�z����GĜ��}.�"G�O�t# #��M�3>�l��:LE���+�:ul&T^kK��^�o��*��8������Z���vɶO9�s71:eKՙz�_1�}�m�������,<zq�ؚ`���N�o�޷EN������M�p�OL�hW�����Gձ�s����1 ���5n`��B+:#Bc�w�;�ׯ:�un�7{��qG�"�e(;�8#��&�J�>��뫂K�E�� ��{�.�m�^�8!f���3MACI�y������[.svC���I�b.jBz�
� �E�x�8p�.k�J�r��鉄��ًEa�X�w�"c	�P�K-��I�OD�N]���q/�@�oK�7����j���6�m��6�\P��`�0`��d��+����/`����k�X�e��tydȑ�1#�C�f����~@�DPҌ����~yٳ�7�o4��sZ|tm������b�W���ؘ-GFi��_h�P���uJ|�a-��RO�I�5���*Ѓjͩ��Vl_s��oP'�Z���Ӽ�f���ke"ɀ�B�I���f�E]��G�	�KGk� d�X-ʠ^�U� �2�aɸ�K0�������Cm���K�P8��]��n0���.�O�����}��m���б�uj(�f�]�ۡ��뛃A�� 96]�����s�l�i~�ه)I=%�mQ��蟧A�{S?*M?�@�Pըp��Z~:��I�{�0B�'���ʗ�Nǲt�>d�1x��؋�����k��4.yN����� �5/��X��,����l�Ү���{�����z+D��
�dų�҅$L��� �"s�"@c��}��Id��ODr�0�By�,�TLE &4!�W�
�D�6�E�×+� ����{�;F�G5��!\��KͶ���ry�e�p`�l�3��@��x����\(a��u��Զa
fd��@�Vm�b�-ؐj< {��1��lE��G����pp��ƌU��b�������W&*�8�4LK70�d��.3_L�Wv�ե���-��{=;VvT@@%�����Z)[ r���zj��R.\.�����a<�Ҩ:>Q%X\tF���Ղ����3��x!t�L�5<rr��	g'Y7���u	�@��+�1|��$��t�Jnè�@�i@�ahU��d��B�@��a*����c�~�9ɼ �Sq������7�p¹���[W#v�L\���VnVH*]/_q���9�#x�T ���x��]w�����w�h�1[t��s���M�K��[��q�`��絆��#q(���V�X������}�������~S}!��t�!�ɠI��+��V��$��RP�,K��&(N�T�Y�LP�
���Pm�"4�v��8f��%��s����2E�ht��C%�i�W�2٧x��E�ǵ1|�s�	Z���W#v4Bz��[:ڜR.�A��"ة���m=�љ�ᮀF_mگ�r�VjUj7*�N7�vl}_+����P<����t*Gd���ݡ4���
ܩs�Ŵ��q1�c���ƪ(t�����MU9��m:�N>�%�� �G�����b�j�6ng�ե��,YK��%Mh�"J�TH��b2/�u�nਪy����z�	�GEF�ߔ`�.�.�2%7cbb�
n�L�7�pNf�b�Uv,Z$���b��n�oL[z�I��6 ���9C �iBѦ����}��$��@�����N�O��_i�7�����j7�n���r4F��  IA�H�I������T��$�u�O�t��h�x]��<w����W;f����fzX� �)��� @ʂH�;)��� ���q����
5�3�o4��C����8���8�o�f�`�����"DK?(�VT����=�S2��N��^��9�8͸��d�$���#�YQ��=e{����(}O¼l���1�O�8GؼL9$ ��ƅ3!U���p~r1�=O�����k~����w���ZM�� #6M
 @{��P�`���L�1�Y �@�8#.T j|����\�\+;h�%�Ox�W�]a�=�DѺcÀ!�� 裁�D�'��Cӽ�q�w�LR?tq ��Q>�<�@�P�vcG��xa��3'-�v��[ V� FAH$�)c�4����֔#[٬5u����Za�[K�*��W�%#l��`���՞]gӋ4�t7�-�|ąf�!�1�0U�ε_E	F!�����s�\��bi�On;�y���� `cÂfD Q �!@)D�e�0dP V| �! �ʽ3#���A�+�Tuf�n�s��t��8j}��6L`��E�)��,EEڄ"�7�f��}�=S��Qؕeu�-ϲ��e�b{v�kV����4�Iˇ�n�"�Dzڊ8��0���;f`&;�< �T�6>�!���ľ��^q1�����$1�麡x��v�B(|g}�!!u��LJ�јpCV�D�2`�j,}9�rb�ND|����2�#�n4��S"I��:0�_�1 }¨��P������EI��`.�?�Pv����P��P�?O����<g��}dB @�(*�m�4��ƽ$��dW�����<#��H������l���Xb����~,�F� ��'�F��>���=�h��&�WRx��%��@Â���D���>���EnH(�����B.j�)�`��&a�2� d�^R'�*�y��S�]R��r�$���)��T����d����<�߯1G�!��ߞ�Y6���E۷��5�@g͂X��mI}���{ZUg������^�Ր|�UDʴT,��L!��T9���^W���=j��<��z;�92�2��5d_�ik�#T���	J+�����z��N���u�"�O����ۡ�����ع�;k+��9�Ђͩ���U��J���Q�f��~w���z��uD�"a
��%&��7s8���g�qc�����M痑��.xn�꼵Q`��TN�U�����v(�N����U�t��Of��U*D[΢�U����51����`UX�&�5�!;�&��������`*\�Q}�|��RR2��f$N�0�e>Zo���)�'f:js&��3�Һ��Ti�p4�f��R�]���4��b�bڭ�Eb��dQu1�Qe���-���l�}�#.��\���Ҿ�vuc���3X���;Fg8;~}k)Z��-C���jd�=�ai�)G[�'��FE�>�.��;1�H�ؤ>f��~s=^��$���P�=�A��4�a�^�#�e� �U�iex�:�4oŽTɑ��-����W�����P+�fh�x��zaE�6=����'�l-����֞�wS����^�{*7���W�~��P�*TQ�l�F�4ȮZ��=L�`3]u7yU=[Nq7p
2��pt϶�	��K$��.�t���)�bs�IV��qZou�\���&Jǈoz~q�����>������8��B0�%����Y(-�/.�_R�������Ш�&�ʛ�������0U5p�A1��,��n	4��j;1z�M^�3j�����9~%�(҇Z'4ڕQ1;��{���X7g�R��Q�@ʌٸ�pBa�nW&���q6�kt&�ժ@�,��7�za�^%%sjͮZ�GY�L��,��6� ����%�m�4�[����a���&��&ұcl]�a`MfN�5��b�j�q4"[�]���LлB�9n��H�lk�7FL���c&�*�X�+��r}�d�(@���]��Z��e�m��n�m.l�v����\[1�KMn�z�n2'��h
3�11�i9���v�S?�1���6�4�Q��Ӛ�}R��i�2"r������(��:j뙘8���"���iJ�1(�M�"�g/z�!X���3<� �ͤ��}���k�g8^�z��@]�r!1��-(,�B�n�t�����u��0�K[��[�M�I�m�+#�C�>sld䥔k)�U�	'�}����ʇ8`T����g���Ce��M����{a��$�=g���8^������r0{ּ�Ee�c9#lgm���AEG��X'�}x�9���%�T�W)W���8E�)���rM��J�pT�!��J�	BP�!�SZ��5;1^*�@�c�.�YS��`��7'����z�*_�w�;-�h�El��b}Ӵ���W�`�J8tx+�ok�è3� 3W�����_Cb�'�T�LNJ��$�&�'��DK0��{/Ȭ�56��"��|�Υ���ߜ����uC`v��CTN/^6��ß��0�2����kM��>�D B
 �	�!:�h�lm
��ĕ�a��Y��G�]t�d�`̘$�`�W}�~�π��`$\H�l��L��n�� �D�C��9Q���/��� b�N��2��{f�C�ӏ7Lw��=ch�r�&�htÂ�{-e·����h�)�x�
�d�R�
Z����ޖ�D��V�lzݱΎ�)�S����u���j�9��V�ꌧ��ͺ����[��R��&0��7N���$`vu���5Wl5��:�?2�󆨵1gj�`��K��f�m�t%ZB�$��wY*G*��λ��P����7���ތ'�p���߳�����H�&G����w�>Znק �ʔ��b�^�A�!�����G6�h��a�90}��׊�ǘ�®�o�W.[a�*f5�.��~˺�R�i(j+��|Q$�m��=��}�1^��� ��L1�Ɗ���&�H���������̳H���0�[S!I�̢��]1Yޝ\�T�C$�ާ�U�w
�w��8���1��c�2�2e��>����w���<��������L�*D�=zg���ݳ�j_������t]���,E`F[�ژ 6s4�c��5-WF��s��ذ��[��{��C�]��3s"KoG��3�{Lx&��#�LY����Y
2�i�}^��`�L�Fd84�NQ�월b�%7
	C3F�1[�j�UY�~��R��q%�ÎjҤLtaG��'��<�ɼ�4E_�1WzOE�l���T7��4dG�ٓXuc���Ř3��'���C�G��&Z	L�i��=��o����Ec�W~C>54�jQ����бI��S����'��ہ�ࢲ��"%͘UK�Kelc�d�Y[s.(�/ ��N{E�͸
�:�9tp�۶UKeR1���]N�	ؽ��u9@nl�v�\�M���DeN]2��� H)�I��4�V�lF�[�Sc��~y�\�������z�HH�	|�����)vΓ��wn7s����u�S�6�p��I�-�8�9D"�.,À��8I�Ƀa�4*;.���Z�k=�S��w�!��(��m٫��	��5r��AN�ًݍ)0U�!tõ�	I�[/��ugD����jlԊ�f}�%�P��B_6Pڃ��H7��u���n�w�|����?m��pL��-g#e��q̼ԷwOF�{}�"FR�R�;�n��F\3^J^c^w���	тO2 e�� ���Ap]q��$��¤e�H[p:�m��,mnM9�T�p�Bh$�T�)���c�u�t\�֝di�w����}u�HV{�����t��+�9���ડ2��Q4�o�2�B�����>������[ӻU�2�M�-���Q��{"��'�1���}�5؈ݱ��H�p@���03��}U�|��-�;"�g�?t�� ���q�bf3Y�7���;��]u,�FV�(��ñ�WCj�y��W}�;�1v�!6�-|uf��&���ϧ�;�6���+�>��1�Z�S�;<}�ۙ�ѱ�%�1]�W��ziL=�y��������Z�)�b��O���<�P�{ة��d4K�ِ:���N�9#B^~�vd(�I(����L"�`���Q˶6DH�nα}�X׍�Fq���D��l91rd�8U��=SqS2Z��of-�B���0�i�!�Q/���I���X�=��cƻSAz�\#=���a�֗nî�k�1w.�wg����SE�@��Y�"���G���5Wu�z��n��U9�G����3GvM-�k���]f:����@aB��y���i�m���ɍOOz�f��k�S>/rl�wV#����4ڥ���2�Y�
�*�SԬ�[����kMtuH��Be����J}�h���i ��a�{xv^|��v�	�ѵ�rLveM��v�����f�<HN�f���2�k��;ڥ�F���ɗ�צc]�nL�_T4T3�>}����89CL$�m�R't�ì;�<��9��K/�	��ڵ}�i{Y�J�:�yG2:o�r��e'u�)[���r����z�v�ݚ�$v�/�݅|M�8X�B�D�L������IS{*����܌����tq�6Y���9z�fe�^��E�JӦb�3�n������W\���ԝ5g�Ū�/��2=����s	(!84�M��q�=�#1�'(ʮ���կ%�J^ٛ�^�c؝t�{�`��Q���Ł� �y�����8z}W��sb��M�S��"@<��
"���@��$o�YGQ�6��+da&3$C&���p�3K	`�֝�[�.3E�&���#T�S���n�ے�r˽�d�
2�K��.2���\,\n�]��5�а�7�uP�fB�h�����>�&tC��^�3<0���m�٢*4n�ZT4\�r�WA��q�闷.�����6VZ�u^��JMu��f���j�V�il�2�SK��5.�i��PѺi�.�k.��+M7mu1.�	�2j�A.��]J;%�����]�gP��S�0�ͷL-l�{�]�I����`�k��K	0����K��ԍ���6|^���:K>�7���l�Mq6ezٞ��S�+�e(�[�-�cT��k��][���� K���S�̗Ci��ٝ�𲝇��>�W6<�}�1��t��=�FrJppˢw�fY���/sAG�8�:C�a����\�ԡQz6a��+���@�1�`6CJn��b�XS�hM�b2+��!�˴�qX6��asو(}ɿ,�GS#aӽ7�Hk�'���y�f8<cU�l|�O��T���Wݭ�~���"aL��b�\�����P�kg���-���#I\��QQ`��-�Tg�C��9{�Z�K�����a�s�D,1�6;��W�X=\��}�"zWn)�IF��+^���ee�S%�"�����
�[C/cd�N�7��׼��#1�����]y��K,8��\�SqU�\�F=B�0�J�iUO[��b�m�8MݕS����ֽ�rPX���y麜o�0'��-�R)5��B;a4�Nym�!��8O�A�c��NnB@�5�b��b;����#V_V]p��0�+�:��B��El��[��Y��wR��i����?:���Ҭa���M�L�D�,r���R?y<�NL6lmh�uf="Ϯ#�w(*�-+y�-��D���%�]�q(��lR2�GHE��k��k^$]��;���밂�M��k'��˄�-� 6��rw+���e�������q{	� `v����{���!F�j��`�b�xLwN�an��2�0��2��3��c��I��ʺc�y q2DW P����^WaI6Lb���㑗sQ]����t]��8�'�T	A���n��u��r�GE��{G��R��L-h���0���m���o�d�@�@�s����O,�8��}�������qc�R|�O�{�����t� ���5Ѱ���ȧ���ߞ����_�,�"��=�?S.���AmV^ꚨ���VW��}ډ��C��|�;/����W��5�ǢG��{����s�e}���Ux]����������ċ����_?>�	��M����0��l���ö�Xָ&�͡�f��kq�;��.~s|�_1�T�@�}y�E��,��qwU��k��gS�v'4��xxj�d��/"�nǼ��Deq���u)1&��:*�"{"�C����-2��&��,�Vߪ� +`�{#�bߖ��!�EE���^�!:��J~F��!��߳���Խ�e �m�o\��{�j��ՙ�u�heL�^=�iC@��	1�u�6}�v����C�1�T
���`�>�5:i�V��2�!�Yq�����1�17Y���ݒ�n�˼�-,37ib1YkV7kKݺ7+j)��h�8H�j�P���c&DT����*@�#�.Z.UC&h�0�ė �(���$.��<�T5U.T<P����?��t��0���C(T�F.�5�ጴLQ�u������Kl<>��~N<�;���8�@����`�,��h(p�I��#A~�vy޾s��j�]��=�덴�E�U�x"�Ͻϕ�pc ^x5�����8(YH�R�g������nV���vwR�1ї�ǣ
�s��0�80�dg+�v�%�\+�,��Jz��"z<�[E�_�q�Z���u��Q����1�>���N���Ɯ�"�;3�앱��'��SR��,U�l�, ���m����Bb�䙛ɭ����.�K	k��!�e��@	�;Y���f��+39��W�'�]��Q��xe��}�ī��쳋�2��~��Ξ����ג�R� ��_ڤ�A@A�"[�����-t���t�1=A��Ѩ��.�	D�������� K~!��@��>=��Ԫr[���[�u��W5hV�֕�ƣ�R���I �%Ǭw������T��ez�pʼ�'�z��HQ�T���>�H
(�L����s�x+��6��X�s����ǉ�AD�ל�P�0KeE׏S8x�%��]�j�y��QZw�mO�4���$��r�z�����ǧ,t��'��A*�*�lh�
��r)�]2z���!��I�@#=S6 [�Ä[K)�[�Nf�ݻ���iBp����A�2�N w�ӛ�^�Vm�RE��m3+�k\Z��@uK�/�����V��׊��V$��n���|�l\���f͍�M�� �Zs-ۂ;M���c���0[m1�tzJYG��黎ƃ�y}�~�E_P�b���7e��}Q��j�}��^�� ��r��*��s[�u2��+�bM ��8L���\�Gt��#��o�*�A�6����>F��	c����:��1�&a�����wY]�<{�\�F8���D�D���������#�VWQy^���L]�h#�b�|'��PftMT��5fFD�K��p�׽�<��EuF\,Y�j}]�xV�:�ͿO�zlb�Y0\4�d��1��η�N�B��s�S9*�ڽU���"�`�Q L��l\�Oϗ�یjb��s�d�����ڌ傫�Ȭ��	�~Ⱃ	��m�[n8w�lfE�,����c5��쎺�)2�i��/�!^���8�mK�v��_-crx��u�+۬�����tY���{���_{��t�H� �!?��L���ąF��'ZM%{WQP�L�VX�O�
�2��TU��cC���������ņ�YHb��*m�FrN��j�J;$\n�����0ʢ�"�-mv�,�QB�e��Ъ ȶ�(�۬V�q�u�eeY�*\�ZZ!=�߃:�MÛ-��(c�ӡ�756��`��e�[v�.�;K�R�Gk�HiY��C3C��7+���٘g%�,��Y]����l�u-����9��5��Ie�,�fsn�\%��M)sVk���86Yu��Kc���͈@u+l��m �ۦ���ڶ"Sa��7)Bݎe����ئlKQn� ,�N̸�pq[-���'�x�![�f��,[U�A�"G"MW5V�c-5��\�X���YVe�`\V��M�i���y��|�;�Z���3��:!V��廸�j{+�����4f}F�z�N����� ��-��n�9'=)j�a��`����h}��RӨ.��#���<&�%E=�G�U��J�ݎo���)��n�����a{��2tϳ.P�tmq�0�3�:�p����0�)��l]QY5��O��
������Y�+l�e@n=�y�Ѯ�)�*r�/��w;������^�]�z��@4��Omӕ�}�������$��! ��d�T� :6<�����m�vG�P���ީ���$-��S��Ԟ1p�iB=�z�=dI�]�����0��O������1�iH-��G��pL��������9M'y��*_^:�W���8��8�`�������j~�9���=�EU�{F�L���md
6z�X��	�.���[s��a]m�:\ĬH��r6�aB��cmL˭�ə�Du��wׇ�o��~O���{�c���lgGL���Id�.9�#���Z�v'�l^����8#���b�v|׮���������@��&I�������Qx�:n���6Ng�N�]8"�GLOb�v�"9�C�G�cu���fVE�*��~ssѸ{r�/^f�$#y��A�@��k2%�t�u]׆Tc��d>��$�����/2SQ�;��o?~Kj�|���*���n	�^�����d)wb�T�,�N'3ջ��vJe�N��h'�m�xv����-O����s��U^����w>ډ��ْ;��s�=L���q����*+*��~�i8�&cJ�Z����@�@�`�:=G�f
>����S� _Z��= �oq�[|�b <��0��{'�*��_;}�ś�3���;n��~�s�r4����\���?��x`�$(e(���G,!vx˶�qZ�#pB;J�lk�.`�jŵ�f&͖AG;��W����ы���מ��L/jT��jQ��M��}K�s������+����S7'(V������H1�;d�Be��Q=Gw��n����Q�Q�U�	�wђ��_pF�8�P���,��/�(5�83���1'�j�z���*���:=a*���z	e�:�.3V�ߗ�+3�^�8��LT�~��E�F�r���[��KN�8~HY�~Pq�1)�q��)w)L���[G��Uk����H��M������!��]���%����F٩�;�-ȕ7�.� ^�05=6#2l�h�12n&��ET!��H���]j'g�̼�R>�Y�f������e�m�=����X|꟫�(��דOz���f�biCnԋ�};�ʧ�֤]ޛ��;��pX�tː7����S���譭������A���xU�����tƵ-��4S�����
�M@i&��f�E��a�u󎩠avι��}C�/w-O�^�
)�m8@����%��z�
��L�ړQN6ڼ�!9�{��F�'�	�����B�Ɔ�؎�RU�R��1��J�`�����ת�<@�=|}Og߾J�g���JH�+�.��N��۫<��mUļ�zȷ�7.9���%�=���$H^�2&�	���(��2gk�_��TT�������/5e�;���yοm���f{s�K�N㜻��.���=ڧy���eP5Y���l.��pXd�d2ߣf�U�H5�G��RPqyj��{�ٙ��$����L��#D�;o�?w�<k��ށ�3wU�8�pn�Z�2g!��$�羗�~�!C@'���]Ųl[�Ei�Ь�1N=��ߡۇ|���}MTH��u5+��H�ǳϴqV(C�UQ�b�w��~7��A��X%���Kd������ӫb�\6��y�\�s��8���N
f�8�P�����Uz����z���}�~E���K
^�N��=�]U�n��d*Ӣ��B��D�xe����X�����l���`#V�u�]cYL)&�$�Y	5�G���ӕ�����yq�]��^��?!Sѷ����3�JfAN��"�O���e{Vs������hA��8��0�z[MWY�z��Y�X�#�$� ��Ъ6�,u����ԓ���� �	��ז.LWx~ױՋ)z/2���0F�-)����Q(�ґ֜�$u��N�T��k���%��M���f�<���LYŖ���#s(C�[�YniҸ�-��˺�hJ�u7V!��UuL�(�p�M����u��uR��-�B�/ӕ����ņ���G���!s�Kɶ.�`��[�T�4���J
�k�.q�w�K��2wf�s�xCi4!0Rqd(��U��ú�Cз/�X�z���p^�Ʊиq����=�{uFz���,��؇��ks ïa�~B`Y�)��[Xhg�U�H�sk^͕��SM�#*�%��Tm�n	��ڍh�Z��Ô"]���+c��1����vܼ�Q$�
ܻ�ie��K����^5g%��9�ԖȦi�`�Z�
��KD�I�{��r6��X ��n��fKg�og��r.�Jk�aJd��f�iW3W[��lf������cSґ�դ.�t���;<�&����m�H�z���j�0�YkFE�T �X��35ѓV��A�r�R�T�B`��;��d��\Ḍ��&�sU�a!2�na@VĤ����m0C����[na+l�9]5h���eit�1�[�$����7ֺOA6��aJ�46�Pf.+R┤Ҷ�����P�Y��+�f`��'�>'���QB�Fı��Xoz��C�g��լ�3����$�E�-y|���h�����pW��8#T�i�:��}�Axy�D���,	L����s��S�M�nmdܭsz��,��K��u��\Y��Hx.�g���*�ٱ���Z�]�{��F�JQ�ޜ��R '��-|ӎ��w�G�����Զ�^�[}*��8���AqӒ�lw@� ◽��`O�e�F?p�`'{g��Tg���� j��a�j1D�7I��M���\+ͯ��bL�)�=c���ZJJY���illuȡqոF'��.O�ڴj�OT{jk��o�CL0�p
~338��zk%W�<g(P/=SRF:?8��*�K��rV|f�Q��p:C�[u؂�3Zr����x���j:ג����z�z��浗j:Y�Y������V"9�6;f��*m���XDl�|3���DwU���/���X6�j��k�q�Gq�R����޽�3w��V�W;۩d`up�����UB���qLn�r0�&A�����-eu���zӮ���@���S��c*����ڧ0��(BۜD�9S���n��ll�D� �~Ys1&���eG�Ɇ��jm��7�&w�ݵ���9��rė�s�9���p�Mt�
�O��@i��Nz��p̺�|}a��]D���K.n�=��,��fd,�Hy�����r��vi�{��ϵ�8��0�j���q�[�:��_d�8򩜩$,��7��aY�~�FǺ�nw�(��
s[��P�I�`��b�kË1����r��5≴|�'������.>w�!��3�7
̲�ݞ�j�-C���g��Β��vz_eWY�{�_�v��oy��1n+��qݨ�`�d�6�.j�ԕ@f�B�-��c~�~����`�c�������~�ܭ�}��{�ﰗ��Iu��y������=�o­L�MoO��
cPY��F 6)��i�1�w~ߛ��MǼ��q�&���/og��U��f�j�n��|`MZ�����~��w�3�e4�ІZ�6H
)�����)ϔOEy#�%v���mnd�ݫ }�mL7�U�aߪ�B�f1��&�R����S�wY�1�A�����s��F��m,3_s�%�2�o�ní����;3E�r�f��X
yZk(�U-��nBF��X�{XND��A%'_Ի����O-�DP������wѓ�Į��ٶGf�u�k�K{v;"�o���j��:9��`(I6o�{,�uV��J�O'Ju�:o����^����|�_S��ݘ���L6sX�-K
}�5:FFsH���R��v�ֱՁu�}2��a�D �e��!�~���v8���u�^���a�B"��$��g\��q��ε�'3<��f�8;0�e
sv��՞�h[��f>�n����k~z�J-��(9J0��)��Y�	tڤغ��mc���h\0Z :|���SFu�U��w7eWK��.RuFda�� [��H�TV.�]�^Q�v5F�ڌ����^�=NN�o��C��2�6.�/�亨�E5��`Lj�{e�r�
rzhk���
�c���ͯc��ɨ���>^��N	�y,�O�r�ow�j*
m"�B.�^���b;c��CQ�t-p��B':Dz3�YY�BS7�j7s��)��%��V�a{���|��$�aٔ�Tm��6Ai�l��;���`��e1�2w{b���r�9q^[+��[��5^��؟ ����:�n��N��{��^�+�>ݱ`Ph����H��h��x�fc{9���=Kհ�����X�^)�'�����7���ƽ�I����@]�0�n����^S�
p�����eE�̤`F��l03�i�ĳb�Ji��-�e���m�m��h��pT �0�o�;�f��=�M�m�ĝ���>�T�o���U��3���+
�q/��ش�tq�0��oޓ�����	d�֊��r��NmFe�{�;���2�~m�@�@��䳴�ܭ��� m_�f�O�]����?+S��O�ͷ�_�DdȠߟ��=&��&x{�e�,��sx�MnB�B�� t+�.�SFb���*�6(�����>�����k���򓕫y���|�2�S��H����a0�E��&7����>^���D��Z���Q(m�k�.��g��u�q<I�7�ݺ6Ɲ�Ӹw�קxW-��ē���n�z��y1V*���	b&M�M�)��nb�7�cu�x���Ф�7�'�c������.�GzH����ۗ�]=3Mp���_w�����E�ʊ�d�@�h��*%?�)��P*���1+iq_�YQi �8�!$�u��O�� t��y�a$�>��	� v�Da 8^�-	�Bm v����$$�i��I!4�'�I H�$$���B��<��W����:�����3� P� ��1����{"�"���n�/�;�<�5ν�븎/����W���(h-;�:�����&eN5������>�L0�DK�M�e~�ǣ��T�#q��y���Y~f�2�G��9�+UPS��ç׿]O@z/�(�M�`��f��H UAO�B~�+q����ړ����	��jC�ʭF}܂�<��oPR��| ��$rr�0���5i�p����@���h{{��2g�x�,������n�(t��%m���pI"=�����Ɠ���H�,�U���}f�y��/���7��Пo� ��VBd	4��+ #$�����2@&RHK	!-�!I$%�	I$>qa# $`	$�B2��HD"I	3�_�L���T>�<uH��XE.N���*%	$��$�'�_6L�_��S�����Zq# ��K��� ��_�; %�}D�lϳ>�	�٪�)B���a��U��^��ŻyB�zwy\��AYr����M�H���J�����y�V����w����u��*h6����6�����A��ZUW���w��\a�}a�I��PE&�)���ꆹ&p�����)D����,a>F��$$�77/�1}��ߑ���0�!!I�GNL�?oD��8	��e+K��?�=��nt��`#0�`g�}���ARI@����rp�X�Ⱝ6
�)�N����8�`H���#����?{�U����&��J9~<�@v;G��p:�N�[Z��U#v*A�Hp3w���
�)'�Y�|围����^FA�v��]��	�(S��^�T͊1����蟟�9'��t��B��O�E��z怑J��KBO-V���1����)B8�%���0mr,4�M0Z�$�X�N&&���*$N�o2�/RcoCb5�ђ� ED�!��q���������@ED�ԕ$�n9�DXI>fm�A@���8�������c���?���)��"X