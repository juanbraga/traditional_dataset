BZh91AY&SYqc�� �_�py����߰����`|�_=޼��7W�,�k[ZѨ$�A��j6�z�@=C�=z� Pj��%Oh��      �O�4�M 4�    )�!
F@42i�=@S@  h$�DF&M�<�MS�G�i4zz�P�6�4H��~��~O�j4�I�i� �eQQ�9 -�Vb �D���"I(n�;��뺟�`H�}TF4���ꇲ꫸Aa"=0�S a3c�V���[9���`�l������� J"0��*��[f*JR��v'����n�ժ��l%e�q}��6-$k���p��2�56�2KvY�nL�d�4(�����ѩ�EA�2RJ�b*��ɗ��Ռ�2�
C-79�wk9W'x�jb��Fq'�.-�ou��k�p�eQ7�����bѴ
���8!*�k�\�s��l�����~��
#$Dd㷋��ߏ-��*�C!)˶���X韁}M�:Z�[�X-��*֛@e3b�M�0\�|R�46��pK8�Nõq0C�'����Ok+�`<��En&6�4��TC�� �	�R�R
,�l��1�)ר"X]�r�<���8iԋshi�ʘ��T�T2K���q�W@�<��69�y�S��%���r�d�@��]�;$��o)�t��[�_=9L�SL
0�z�
�$�7:�`�
u��nҞ� 倦b��<�-�O�1N�Jxv��A�1�^���'}�h��*f�8)D1"�0���GopoQ�'�x�VO(3$ܘ�1�a/W�����T���ƒǎ���t�*kb%�^��ʻU\�+�.��e�9�M�!"T�nMe�K��]bIY�ؠf�s4�[le��f�B������s�6�#����d4�s����I��Ի,�.Ҫ�;��]Ƿ�_7<�K���q�W��(DȖ�v�T�@�1S�9v��#d��*����ĵ��T�)/IZIYL�M�4`�jI �%���h�κP�T!UR�0b�@�Rb���.�R�22��Z�9�EaL`ʲ��K싾��h����4<됃�7E�����e�@_�w�%���^\r#Z+�#z-��oL��\2�!���,q��t�$�'���9���Y* �r����p5�����^#���Q$Q���Z~�#�l�kM�wS�0\�R�oݠ��
�r?a��O�R���y�?.���.3�%� �!�%��pn�x���4C�̦�s���D��$�u�S���j�]ϙ"�� �=���J�y�Y'�.P�*�T�AS�ke	,V�Lƒ/+ޖ(�y�_�=FF���d�(e�;����9�/	[�A�+!>��yz�Z)�-�*�+�"��4/;�4��0;v05�V%�F��t&I�O��������3M��z7tM�v�*r!� r�@}��t�9MIY�3&u3���z�J}��Y=q9&�5HG�r8���:�ԜP�2S��Q�n3}�%`c�jA�Dz�Ѧ͌��$��MqeqR��@&�I5�ә0��ȶؐxI%Ψ�
P��;)I���2	ٔ��q�Yd����J`!s��;TG��P�x��&W4m2c@p�p��[�Q�k��=��%(ߟw" <��@�H9�S�~��(�ӻ��]jB��:/1��F��eF��/�7t�6(h:�S-M���$�F{�U'@)Og#��baХ�c��_�@��'*���H�E��&˂�L1�(����I������\��e)W]]5�fJM��\�P�d�5@�c�|Y=҉=�}$ ����-�+�9M��:�k29�Q���ݨc9�&@rX����]��BAŎj�