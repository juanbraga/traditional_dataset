BZh91AY&SY�'�� 3߀Px����߰����P�vӸ6j�Ws�&�4L��=O&�jz�0�b�ѧ�D	S&�{SHA��1 ��  ��%=&�d~���I��M �@�4ɡ�	���dɓ#	�i�F& �"S��)�!�=@ 2 �"�bZ"H.Oaп�;��#!���.� �0��85�`��4�v�R�QN��DK~˦����g{4a�5�-ԃĐ��h�wR"QJ	�<�.o�d�%	��E�:&����fL�ٔ��+��3N��8��S2�5���D���;@�1�I�HT�1��դa��8[X���5�+��ܩ\��X�L��^\�����6���z�2S�Q��b�gTRl�>K)���F�v�A���,��K�ԃ�4��Z���h{F��[�w���K��X����ڹ vo�U%�l��t>��"d9�^Z�r��m���|�NV����?ۤ4	�y����}f6Tq����ެ�f��=����(�d����S\]�Y�Z$Kܙ��y&l��b�/>�kcv���1(�pXt���g2�U����~̘ª3_vy���ɡZu�8F�S�c���0S=�8P�
3��Q�&D�}��}��yw*g�K��׮.�Rqׅ�|�x{���X�{ӕ��ɆK+̤/8}�'p�~�%�׼����yM�*�(�m��⾦Қ�i�\��K;���*��A��!\u��K��S��cR�������/�<A(�Գ�	0���v����K�"N>P�&1�
,�n*ZA�E�%��B������5ܵLj ,+(*���Ϣ^���Nz�]դl8���I��m��}t���S%��*�C�4 vF_P�YNP��2�*Dbq8v�(
E��p��/�9�BiK��u��2�[$���7�Ŋ�,ݤ�{q��QV@Q����-ҁ�n4�qeMY�YAB4Z�O�U\~��=+�0��O!VUk�Y}�Zo�̶�(K�lNfA�ɐcG����ܑN$ ��s�