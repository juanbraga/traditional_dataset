BZh91AY&SY1�Us �%߀py���������`d� �	U{e*��h�     1�� �m��5�j��Ӑ��t
��@�B�Uf4U 
� �&ٓ@-,�B��VmJ��U -�����(�4��ʥD����U, 3I*�fb�S)D�fII�) � Se$�2ԊR�ePfi
+-$$��*[� �TE?	USF�z &�@�h LMS��R��� &C@��4��a4�C �a&&CL� �Ѫ��D�� `�L�d$��@L��'��M1���'��4h&�MD�24�Sɦ�)��4���=COI�Gl����G�@l�笐�H0&`HI	* !��2�@�G�O�4��BHI 2����´O��@�C�$)��L2�H@���������x����Y!�H���$H ��H�H�U	9d��BAH�� 
 L�����HR-�� P�)�X�I"��
�Ba RB�Y$ �!h@���s��'�QA�q옞wo~��uxf(�5���]�U��tPu�ʛ���˒"�D�\�)���Շ$��Q7��/@KT\�W �&j���ٺy%�0��bi��6ӌ��إ(�/(��٪�Yuq�� �Rw��:�2.n0ؘN(a��&��c�+˲ZS&�.�(f0@Fqk.^�&��46��Sx~�NDW�Ħ���'"�$Q��J��"�wF);�p0�YQG*��B��'���𜟩�-2rA�R��b H �S�/�!:����iE��1"�fL�y��6�En��ٳ[�k�D�;5�
ƶ�NXb��1Y�Ta!������Ně�n,hcLKGq5Z�Ԫ6�A�h�Ybc~�Ff`/�
̸��f��,��)��@�E���S�g N J�3��Ok�D����M����/���TM��Y*���X�Q��@�Q�1m^��h�9%ź�qj�X�Aʕ$8�TF;�܄T$�r�*X�P2.T�5��VI�J˶M�ʱ.N0��T�����X%�Io�Jn��ڍ���|]�;�EAn�*̺q0`\9E��6�.��̹���6&���:����Y.t��3rf�DB?LR�pp��B���؛s�&1M9��$9��!4'I����L
w��Ȧ��j�oV�7F3E`��-!i$6ÖH,!��j�ZCiXR�!�T���8I9`He!LRm�?E�^��Q��b˓t�d�Z��
tA�p�&U4��w9NX�&��(8�����	��'��[iڵA�[��^��Qve!!I�Vb�@�e�pC]D���c�A����FSȧtLayd����Y����c��I����o�wL�Ci;[xYۙ��ۄ��w0��#�%��ꄼqn�A�,Y��b7V���I��Ŝ�;P�mR�5�'R�`���]1�LĘj�(3V���®K�8Y/�EL!�;�V��ظ 8ݗ�^H��qS	��Q5Jud�k2R�NAS��MVSH���@�oE:Ŧ��;)��.�Ś�����bV@��p��� ��q6�S&)��I�R���\�d#h�$� ���[gE��?�~g�
�N�!֯F;q�C��Y��°8��Z3A��y�_*�UE]���-��� ��ۥ�n�\۬frĖ̴ei�	v V�֙{�F��B��M��#M��&i�j�q��ܳ3��OJ��j�\e	k���������1b&�[-Ѓ���eI�5cÍ�3InQ�l���q���c6�XRn�K�m�Ͱ[Ƭ�I�8�	u���]`�D�Z��-h�]͔@��J����Sk� m3j�ش�[�u��u5s-Ë��"��Y����n5hK�uHY�#���P���"��m����F�e��-v�b��J�v`li��왕��D+uM6�^m���Z׋�J91�n.�F��P)�ىkk��k�F�qt���J[2b���KMs�b֜e�6�Ú;`�7�k��g�ͳkV;=K˴�Bn�[�,��Bkv�2j`��1�i�6��f�KUh+vv�il�in�c-����,��ݮ��(5�t- j#\�b6V&��ݡi���jٺ�%�)]rh�,�`���]4\��%�2k�+u����$�s�/0��L�X9lbk�f����*陝�U��tcK���]=���Kv` �F�]v���<�<���ʋ1�^+�mj�^:ٲ��6�j0|<���΍e9uH�X�F����jL[mY�k����I���PZ�fx0�@8!z�P��Ax��Q1��iʆL�C�H��h�cu��]�ͣB첶]0ཫm�+��.���k`�,�k�S5��JYYlXK0���]f�s��$L��.�e��닛��:鮊Ylm��X�bMp�6�́m��0 K]Q�)�L��z�M�%l��������Q����]��!H ��a� @ ����$3� �>�p ��=��HHAd���d�RCΐ"� Z:d))w$�a ��� \�i	S =,$<!��2�$��!� i�m a��E�	l�
@�@�� i�(�!���)0ɤ$�^*����	#��
i��
dʭԽ^�SUI�T��Ɍѧ��8�,���8@�c����6|'�O^{��$�5�5��DC���W���L��
O7����^I��!�Q à�d�51'��@�: ̓N  �X\T���#S��5$������
i�C�RZe�?���~��~_�$���a_4�����'����㼞���x C��o�T�~(|��*cѾ��MNG�ioCn�!s��^ѺQ[u	��Ƭ�� `�u͎-͛���@YI��遶�k)�j)��ל��ؽ�v����fF]�blm��\���m��li���I�ؖۄ��l�L��7��.�ҽ�)u�P��7i���56�%2�֛�9�L!s��%�Į�6����b�n�]萁 �]���ym�M��ڜis����3,۪�#[�in�ŋԴ�RU_�ݒ�B,�e�) ,(Z�6�±(,Xm�hp��,�"�IB\k��e�W	C�)��P�J��P�ʋl��+ULFf���Ŏ9��U�F"*2/�ҦR�p���"sί�
1TB�����(��4��F%�[���R*����P�)J��E4�(�`��4��7t[IJ*"Ҕ�Z�� t��5)8iW�j�t�a
b��Z��b�5��9�|��:��.,� ��� B�l�$ �<��,��<>��纰��Zc�m�8_{0�'�ϧ�_s���_&��UEz����R:���4����C�.&EIm�i���mE2�T����;s���0���
�iL�b14WU�昙�̘͔U*��DD6n����"Ȉ�q
 �Qvch��d��i6�1'����z���nf4[�g	LQ��VUQ�4�R��U�UCCiz�7�T"UP���5��)Si��s��'I:�z���3zr2�v����3c'gl�EJ��}�N�N'����^��'��{���!|�ȩ�=\��wopΈ" Fn�U@Da�ueLWM�VYf는�p�X��m[�jL2�]dp��3�� �"7��I��j�$EW��E�1	1I�K	�~��M�ϯ[ȓ�  �� �a�#r��3�f��Ñ�x9�T��XZ�F:޵g��w4Y<T������}!��0 C�1Dc�"���L
��`4Y8x�Ny�t�öE�7cTP�]uK	T�� �01{e|��KJB�M#z����z�����q��l�����c1L���蘎�$��* \�%���[菬O[�J�YN'�{��ю�"u#��X�EM�f»#䌤�`�u+�9s*�e[X�nm��f,�L]��pj3Wm���'���[�/�7@����`�egT��"�o�����l�p"��îȨ�H�Dac�!�f
g�r3�+T2a��� ��L��Gɟ���|� $LS�U�0�*B�;&��UʑÕ�Xn�@�*?�4��C�
�ɫ�"��J��Y1�-�ε|�矑x1��i$!η\_�(�]�%��faD֪���`��p2\{<�%����ɢ�����`w��& Q?W)0"'T���[T�~�(̟���1C��)�	"@e�x"��I�#�-L1GUZ��Dt���`��M�r"U�LF�&��bc;�˽1�|\}k*�,���B0�pʉ��k%��~BI&q�cBp��Ɯ����L��͗iKUӔ��޺Š�� �l,c[{�����·T��`F�gW�0���w0�+��u&���m��I��<5���S }ѽR'�� �Q�	��*6����Au�^��d���_uv�lR�.��DH����,��0���-��bq��z_N�g�⩀ 14�zbEJ���d0&L�D&�MN�E^��LM��]d�@
����T\�tw��k�y2:�	&J#�(�܊��I�,�
U�j���I4R�on����0dc�,��-��x�nf1N��Fˤ��'8�7�7�[jsP�o^�E��]��p�bL6�+q9yĨ A<#Rqzwp/�� ��$�8+���|'&����a0� �`���u��	8Jd���t��7)��]5�d9i��rl�N3\3T�I���#�d�<�j��}8.RMi�&���R�ĵ�
-���7�z�`F�TL�	u�J���C�5� �1\\0��&ڊr)���ñQ��S��s��}@�R� �J<���5۫"�&��p��}��=�?+�zv}"����X�NCԇ���j �$i��p�q3�kr�䈜��x/#L'.�!�eh[Z��P�ٖ��T;���Q���R��Zͩ�ohʒ�H�9��
�tN�v����<�R�iX�&��n��ֳ;pVݽ�o��R��4�ꂵ�sxg1P�����[b# |��b�[�|t����p��ï#<bJ��@��~����������G�P�	�2}iď�`��hP�Ƅ�H@���<���u">�1}���AԆ���B�"8�%]n��DS��c�c� @�Fb�DX�gBڏ��{g'�1d�����z�y֊���I*8�pa���gK�� ��@@��g�5��V���{�ϲKoD�ϟQ �)E��U����� ��Lؙ��_�1�\S���O�O������y��F��B	1�1R~�6Gĝ>�=�I������o�7��b����9]dO�����Kl�5�{��Ԕh@�>`CG����> <[��L��PJR��m��m�Sd�2R �a��`��QnnN��65+2(
RԭQ��W.�� #��#�>��1'W�ŏ	\~���z�p����g�DQ?1��"��C�#��`j=�E���eQ� E�#��2 �<O�&�>Fz��+J���͈�0"��&�"	?p� �i���* 
�L��䎈�&� K? �")�kn���J�)	��S�Y�~&��|�x��)�V~f;��i�op@�"l�/�fcg���/.rU�`���<"�W��L��5D�Cq��;��ؘ̺�v�⠐�%ez���.��	,�e�w�(�,�PI_� V���	xק 4�Q�p��wӂ�v��^�C�_t�v�ȥ�	�i��*G��:;�s���U�2Pԧ3U�Y,�n�ޚ�C҅�QAԕ.��PR�6a��M����9��\�O��xb7��,���Kl	�F��v���$�]����`
%3�
�hvw^��G;�>��4=8q��7v�n��'�sm`�Ξ���8 a��ھm��ө̬��R�ub�����+��6-���P�`���Ukcg(����s�Z�|���KfL��ԮT�z|��֚��޼l��=�v�	Xʑ�.	aZ�]�9��5���p��M����"�M�M)Y�5��Ź��R��
�ꍽ�լZ���n�s�ȪQ�-�B �b�x��Tۦ>K�G}����s�[�d��O�^�8ɋ��#6I0�i�f�������������P���ĝ���|X�,�}�U3�q�jhx��9���ы����j'����]2�����Pt�����yqb<,���A Zo�;-P8Z���N׽�W�ZXz��ώ-P<��0tz�=���A�q��*���$����lU7q����l�CW�w��pV���a����4YI8���)Oj|�ޘ��^M�~�`ػ�H�j�uM����f	79n_���̺����L���x	B�� ��e�!���ffw�W��V�G���j4H7ʪ�1�_�{�0_��\��7yJ>��ϲ+�\�}G�l��ñ/�a�1Oʌ���or�0j�|�2�A���~�	�eY�ǽ����]&[/���7�t�)�H�R���7#U஧}�����$tQ	�͝��*f��,4�d�U)��.�"�n�"k..A[Tl�S�9&��f�ڣW�wKWnTK;:�4Z�ak¥ݫ$am>��lX!Г�ָ�0�m�iNm�a�E�Ej��ɡ�P�U�Jp�Al�P��sjl]I�l��`W"�at�PU\;2�إ�k"�LT����4�iRq��H�f�\�L�ss@�f�Ц��di�]��Бط6�*h��*P��ɲ���-�[�nͫa�C2��f4�t-��B��cYh���A��(Ab��r:к����kj���0���?G��]=�L[�t[���y]l؆�Kuz�3jg]�31E��\�FWaV~�����~��G����'�*k-���P���b�ܳ|��1�U�~Ex/���ۘ/sƅp���4�G�l���(�� ]���<�pi��OW-UP���Uдp��B�P T����Cy�	�Wr��C�hHy�:=�s�Ui�L�r,�'/�ȪYp�z�q����b���װ�":�Z�.�K��l�M�0�hxTܗ"_�l�����h۶,�����m̦����2�)Ǎ��l
�"�p��5�{6=BYXM�\�jy*�F��0��Y)ő����jAw^�p �À$\Uؽ�QOp�b<�|7 ��^T�6 O]Mg�$#?7���7k#%�J)���V���@~r���|���/P�9��4͘�1IQ1��#-q�AH��٭��ޤ����{���=��g��̭�uy��1�ތ~��e��!��G�筛�߹e�QCs[RR���z�/���C�ֺh:��s}um�l$َ�-����˭�iktbݚc���[s3���6��A��c�p:��b�����{PMo]9� ��]2�U�M�I��j[����qsu���dhIvMW���خȹv��/�Ȣ\B'�v)����_U�nW�w��q�5[۔�Q��ejS�8v!N����L�z�l�g���K=�='�*���|���7 EO���q�̻ ��d�_������mL�/}ςM�	"�-겶�'��nLUI򫪳c�6�,q,������w�$D��Ss�]n*�#2�d�~S?^�eL5�2���gc.�B>�������������g��n&T���UL�O�w�~��] u,P�gTn�[�)��<h��q��;���N���mB��9/_���hg��en9��/Mt�$Cޣ$�:��
�N㴶m�8H����ERS�m)���N�o+e��~ ��`��^�2k�L��&'j2D�MGm���[�ӣX�O�7�!�J�R�瀀�߼p!M��`0�2��!����;�]{D�kH;���Kn[E�6snL�l��=B�};�|'#�����ռ�)C�ݺ��9퍲�5��,�ؗ^b��\�{���{�'��oay��|��)�-����y�������c4}B�{�#א�nLw�Q�X>����9����wD��&��g�$O�����|4��:����U��@MM�ީg/�S��DL�������+Q�b<��>�3NM�0�4ys3��m{cw�g1N�5�N�	ve���2�ĞF[y��l���6*-����%k��UA���%���2���'�bDIXq��]\�d0�&�0Ӷ*�����-��=D}b��^������9�70}͚G7�ִf��_u?n��m�NI�R�579�vSI�v��zv/Nj����`�Բ �md)������c3=j�񜒝k�\�zR�ןdg�}� 2/���*�*��v� (,��7[ಡ}�%^�N����b�����Y����W����Et���9��k�HJN�v�G���V,��K��X�v��3a.P��-�U5����p%��.���T�MVl���2���] ���s���wo��k�,�'Z���<��ztb�V4Y��o�\uW����C�~���Pױiˉ�("�$ӱ^�!AP���+V'b\�9���Û��G��^����� �������)���J�7��x��f�Ώz�I�]��ὑAT��i���}"���D/0	-��i���o�S>~�*�z�oJǾ�Q�4=G������䴐�أT��{ >��Z������x�9<��E�{��瓷O�����ob��O=}� 6 ŹX�k�jjGF�U/N�1�'�.�&����rc^��WF�_��Ѭ�%6��)����Y�jsl��G/l����|d�v1�E2\aZ��^������0=A�����F��܃�gb�x���_��A]�4,��X0uǣ��\o鉔��q� P�����x���/��{Æ ��^�:��*6��*д�F`��2���چ�A��K�f���0�*��F��1��Ͻ�w�>���s׬�܊>ͫ���=����'e˂ό^�U��OM
ɟc�Y�GzW��	�a�@;g&|gkv��r�2�� ��{-?�T	��c	����������T�K���j��}�;�<b{S�@����Un   L�Vc����Mt?u�:���*	go�?G�<v������6F珅yE�����F7��2w����M@��:�~�>+�).&EP��"�Ջ��fo2�4�^�%jk�<=�5��]�C�3�|�;�p�lz�+�xqͰl{l#U��"�7��:n(�����2�h��>*!��P�Q�x���/O�>=�0���=۷���nAG��4��i/�q·Ĳ�:��p�x�ϢG����f&yj��2\Ēj�����O�$����~OߤX���H|Y��&\�����,
W+-���'K�%�\J��2�f�5'gv�㓆eN�715(]��we�!��
w��v���TYj�:�a�&���ͫ,ɸ�R��#�,���}}|<A��m�aШ3Km�ݲ]k�0Y�Rb��&�Ƅ�!̤�1m�H�ʗ��k��hԌWm�j-�Mxqhk�]��S\\�ʪ��1
ʶ-M���*%5)������ck*�P�hÍ�1�j��Ve�q61bG���4#�	Zl������"i���f A?S;�����y"��;BĀ�Y�����A���n�Ѽj��v��I�`��ۭi.���S�1����SokA����jRV���܋�~�i��;����[;;V2eG�H�����m��I�l�i�����H�ZP]��¨# ��=NnӗY1�_e���˞��F�o�2��{���Q٦��U5� �W���D/��v��xG���8����.���6&�+
|��*��8��]�h�ĸ�P�f����5C�Ǥ��C5ز��9|zB�#���e�]��>�C�2���i�K��6�;��| ����+��}#]u����E��38���]�djԸ� s��*:g��D��rQ����a��FG�'Hi��_�%#`���K�'����)1�{o�iTz�E�{()�3$��o.�����*��B+��|�d}��׻�����c�գZ��,�ʱ�3�qK�7R�c7(�2���K��1w1���}������~\T��#S�CΣ��
��}��e��d�9ъZ�H����K�t�ֺ�/˞R�1xG���{Lq-�B��AŜY��e���-��wY�慀ڞ�&]�PR��8:68�F��k�\����]�˳�Ȍ*S��S�J��s�g���=�'�)�T�%���ps;�Y�)��lem�K��5]������cMo��
�����Yz:)��T���z���'��(I�*�8"HCZaE�аϯ0"������Q��Ty��wϦ�d����-OǞ�rۣ&K�
�iz"�&=I�{bE�~O�d0 ̫�uT���T��> '�L�e�݆�������EsE
{��Y�#wҥm��oՓ�}�W~�U�8�/�l��	��*_[��Zr�`���3�޴��E�@�f�*�H�]�,͌1khi]�.iQ`)�I$�`���U��ب��Cy���yv�f��Z
���H^y1��X��k�F󽹞�)k>[�s��vv�*P�wd��ڻǇ���V�S��w
Y�Q�V#��Jy#G8���z|���o�Ǡ2����"��߫��
m���*œ��J�,�)KL�_H*E��n*�^W'��"C�;�k�=dq���d�!x-�m��a&A���_�1����b��[s��������c�c�>��ׂ_�u��Z�#꽻�Il�V�7E�i�sjr�ԛ��W�)�U3{��˔�jjZ�(#�w� �H`a��/<<^8���I;#���2sY��9�:��E��p6�4����U��6���}�*��9&:7d�����پ��d�l���&�
��tv�	���U燼w{Љw��HB�˥�ב}����l{�#mz�3[�����8��qS�J������56X�Aq3ˍ.��%du:�˧j͕���$�M�����+mC�=5]ѻ�baOd�*���İwPy.��Ē�z����EL1�MV[�̅�ϸ�5���=~��aObLt"�"�h���v͆���u��bY�B��b�
��5ֱ����~~o:{�>�Ib�����,=�q�鸛���X�E��B)rt���F��e׳�]Ix��7d^��hH���sB�YZ�d-����q�s��26��NW8�$T�H�Sf0�w�ظU?�غ�{o{Q��=��=;��������l�P�[�2X�P}3pB���~��#V��ɡ�����9�<��Q�B}V��rEk�U0^�y�����Y�����X3�Fל�e�0�'K��M��B�M�+L��E�]! ƽk��x�v�U���ݰI��1r\�2*=߲��s�k1��Mx����ІP���e�*�
Wu�qպ�MW��ɪz�G�h�5{�>�����ٙLc�h���k�?o�Җ�4�)ĺ���J�Cp��tR��BJ�`� h'#���<G�Eu���䔌p�+��35��\lX�O��?5��bn{���={�=USy�5U��s�?MR�n��<L�+�J�͍�Pseփo����Y,cZ�g @$�z��+�E��ALsN�
\nu�Sti��F(��r:Î'�_������0�3Mk�yJ(ez�ea�	�J��ӷ�7�x]�~uݝ��t��_Q�=q���ȿO�#��v�_.�=��r!��O_V�\�hJ{Ҕ�u��wL$#>,8M5
��Rdi�TdQ��!]��l�뜺���{|3��l��qmF�ݍ������4�7m�+�B[�ժMWY�fH<��݆`"O�R��{=P���|q:O���ʅ�f���r�я�]�ᜍ\�󚥭��7�R��ŘS�0v��q�Ȟ���]4�W�����WVB���2�'����-Q���Lё�1L�A�9Hm8���QO6໑�P����1;N=�!��8ӆ�Ϧ�7_l�6hՎ�V7\ΤE���q���
�{Sfw2��YRa�KM��L�e�'g�����������)�`Zh�n*2�݇�5-��2�X�khDؖ����I���5J���z�A�[��V�m��Ьq5�#2���s�]���4nЖmT(5�a���pY�f�:���qmk�%��k�K�/f���ղ�X� 9lͪ���B1�ֶ�t��L�����[<��k\-��v۫K��0��K+wk�nmF����1�XdM��� ��-i"�v��GU��ى*�-�c%���鶊��0A�mez��ڼ�@�U�o)�Txr	��m�~��5x]�;kze�"�tM��P�:��'���c������rƪ�ܾ���w�*�q
���py(��8��Q0�U�.e4�p�t�Rk�9ʽ�(��a( :if՟e�[���{p��6�ǳ�S{�6��A��Q6��JI�/.]Aޙ��Њ-�J!2&��|�=�y�����'��tO����J�����p�`-����K�Eׯկ�;^���[p�JzCs�(�6f΁)�q��.����	��I����Ȟ�c��U�F�軬�<F_>��^j���Q���2��/$�z>
�46�w�>]3�E�̘VE�	�`	���l5�!i�4��YY��fU�Պ"J�غ��x���'x��(��zz�A����]�U��]1k���cC�ތ�>��ӽqsok�c����ۡ]jzk@��0�6�Js�=�M������;�������E:ݗ���S'f�#�n�r��I�uG)]������C�~㋊3h�Y�j��AGa�SH�[{�Ib4av�0h�gI��7��Jd�hx�0�a]XnWf�������E��W�Ʊ���_T���u ֪sG0!�0
�PM�q�6B���nR��䉒�i�~����-�j[��U�o�^�ΰw��y
�o��E-*p�
f���Ř�ޔ�+�%Y)\�[陰�S*�����K���7���<#׾���Nk���\�Υ�6#����&0c��Oyt��>������������a���dƴY�k0a#����m�k�3�ͳ�6啊\�ZFfշ/���_�_���^\� ��)Gyp�.��l��K����'�me��d7�B�f�f��f`�t�G�t{JE4�A ��4Y��r|re�Z7�{-̕A^�{�p*�L���o1p�p���b@���gN���U���Vs?qR��R�B)�N{H�T=y���d�i�҄�����V�h�Nێ׹R�VdYs�0>M�o[l�
Gp̄	vʽ�ƅ3Z+l��K��墄4ã����#���U�U�n�m���:c.(�٘�̄Jťd�hz
��ɍc\ӱ!�]sl5U��K��ٍ�83i=��`�e)p]O�Bj�9�*�_ռ���p�lCi��޺|�fq��wMB�;���i��Y���:�������{��������FǇ<Ƞr�3)�8��y4L"8�fqͽ���}r�&��"^�Ǝ/a��M�! �a� @뺷��R�m�eW�9�y����7�!���z!�M���,�KdՔ��֕��M�]	n�W8�m�\�?3.@0�$��˴4]����Y�&ƫa�o%g�(�t�^�p�y98��$�Y�R����\%[ջP�Zm�é�b�=){�}�2�s���R��B�o�	o/��z�m���3c�k��r�;�y�w�پ��������+�|=W�F���C�H���nf:6�=[�g��i��G4��ٔ�����f[�3Ќ�Նno9���������}��Pr���ؚsP^�nw�$�$�%(�R~m��uq�Ѳ��7 R
G�.U�}>6f3ri�س�Wt)|�|�b1)��_r�x؍���;=�R�D�!�Ѓ����z�l�4���_e�*���W����Kw<����\N���̯��$�>�������۟'�_<t����a��\@�C^C�������Y����6	p0�j� �>b�xT�����h�[3�{ʵx��9���� ��?,�U���5��pE-ᗺ'EһW'ޮ�h�l�����-�Fv$����/(_�^�M]t�xZ�R��o�`���gl�QX�m��t�\��+yl�u�#�uã�N)��hǟ�v�(%!��X�lϗ��������|`GWF�Q�v"0an��,P4��N��	0��a��OΚ�Ƌ��~̼��W0�CJ � �W�&2{Db�~ĵR�Ë��gZ�@ cl���Z;Ef��y=Jrmd5:{r{����V�Z(Œk{%2�4Rw`v�wDQ����t�Z^����'ӗ�[��Cs��y�5>l�y�厶��J�����jf�"Ε��b�u���fق�f{1�c��7���1���Pfܡ8����ŗ8	Q���Of�6��lI���Q�~ܤF���c�ͧP��b��-i�F�$2��$������fnJ�j���[p���!|�0� �0�붍e�f��au,f�c�..�[ƶh4m�6��5��4��.�L1�F�i�T�0��0�l�����\%%�-l�^"ِ���`����l��6��H��#�����Q҉WkfC[�aXV�#�yո[��lZƺ�ԇT�m!fA������16O����k 
�h��CJ6c[�]*�je��l6+-�U&�`�_h[�R��|�����Ez~�plwb��z�=���wʽ<��%3������)�u�ЏC�E<�':��D��!@JN��路�d�R����Z�GK���B��"э�Q�<�K���jhK�n��@���Ż�m�lTW��K��P*�
PT�R�H�5E��}ٷpD���m���q�]y{j���[ЫU�Qe=ޘ�4U��B�fN��)��s	�XM����[������֕kU
*�*�q�XVK�1���~��v���*�LwJjlN}���8�ڪܙ���p���`�����.z}�M��Ч>��6�:�#�Y�}Ւ��COA�~1�}~�Y�ü余Q��z�X���Jgb���I�����IC-����Š[k�Қ¨���d����Sj7wϯ�z4i*f���xb���⽖�	欹GI.V�p�\���֌��e$`	�9E�%���^cȢ�M��m��5��.���j��h�wU�컱+A	)TU�^���[4��`���Wu�{޺��d?S��`N���pQ5²U���s��c�&��%�ɓɉ���tl;�����R�LYs��+i�J3N�Q��/7��:<=%��TJ�]vU�,��(���-�^�zЫ��,n^�{C�ڏ�<��Ո��oT���oY~�{�Wۦ���T^�
7���z��S:��F� h�Ch��p���G�j�tȹc��įe<IP�(W0�f���������=v�玫9�M��a�G(�Qmٻ<�߂��0���9��P�U��q�qmx�k{#Z!����������U�y�8z\j���=}�f}t�**�Rc�-�sT��O���K��^�M���񂂤I%"s^��|�G���"�>ƅ�)���q�i�Zg1ir��LOV;ؼ��6A�۾E[FGv�WԺE���g�ex�	A��;�S[v�ۅ�y�t��{(�թI����yS��Ň��?$o`�ɹ��dhZ.�No6�]UѪ�*h9sB��'V��ր�MM*SR�V(V�3e6��Ǵ�8ʽC�D�36bB�ʝ9�D�y!aT�l˄F7uV�����ñ�e4��T2��T�J�~��iVک̈́�� �v�0�:��&c��z|�H�����.eK�~͢�,������&r����l �͛�e=;��=$;��eI���]�ˍ�7o��yQ������#�va���AH �\K{�h:��1��[ٶ�+9⻤p�B>>w�G
ܷ2v�E袕����<iG�6݊:F�?�Av6����A0�ɠ�.���L�5��k�hns�Q������ l��_��Uf0w̏m+�[��O��\N�o}�5��xu�!&iMY�� 4?�M[U�9��ɕ*��c\K�����QѹN樷z}�r^�ũK�_d���e5�7wJ����G���Y"���λ��g����z<��p�~U�7,�{d��tmn�u��\�g�30�7�r:=��Ҙ�o#$��F	N	)�S�#
Oc�v�z�}���^��:�+t�����=�k�Wݣ��W=��`��l���ޝUz�I�«g�,˜�ˍrD��?(-�K�fS}�U�\�C�n��}UU@j��t{�S����\4ZO/�ʜ^�W���Rb�͹�<��71*|}i��&��ԄZ髡v,HB�vբ`�[
��r���l�Rm��I^���[7\�V}�9o�8nW�n���I`��ݍ��F���='\��Wh=ƛw�G�E~���.&�-�Q�(�c6��΍έ
.�6B]��+��Y����W��}�qz=Lz��T\�����c�d���JHL!h��"�q<�o1�&cb�)ހ��t`����t�25�X@M��f�2��}�(,��Իq�2+F"c��-�	�cs7j��0�=h������d+�t��x�m��.�;ik.�Z����1R�LS�����<2u�����"�M��
d�RB�L��Bݬ�o	���J�(���B*�����Z9�1ӓ2Xy9]��eE�C9�G�����Ԉ�����"��U�$��B|�Hw�7w�$J r�{�%R	�/�� $��p�������8`Da��@:�$�X@��@$)	ބ	62CE2�XXQ!�J�u$�MI
AA �w!%���ʜ����P���p�|�}"H"���;S��ׇ��u�	墎F����{����s�r�<#}��K���%x�������^�7o�f}��\f,����S�ZI�À���<l�%C<<����HƢ���H�BIZ�z��z�)ۗC%�=|� A�1�I!$������''���g�<���O�L<)�dzR �N�쾕�1�5(�G�==����$$�;��}I�~Z�����>�	�T�~'��A�%�Ώ��S��<�RNpJ�޻�����,b��'�9�Ĭ9�����?[v��w��4���L���]$҉��?�r��T�	)�4s�Iyt����ˢ�p�H� ����ۤ�&l)���.2I6i@�����E�T�BDw"�a7��T�Y���ź��Wec[�UoX�l��w}����� 
(�����I$�� J� ���.�%@��F I�@�I��	$�H2@������.�G{���6(��S@�}�Gl�@Hf�T7�5��D8&�YGt�I?����(|S��3�Y��N�>�����䢄�F|�_������!$��2��\�¦:��X/|{a ��qE?i��d�׆b0X�BC01�H�? i܀�(���?�{��HI �X`ə2��'N@f�{�7�b�i��h�bpbW�$�H}��@���쟀J����>��5w1ȕ$;˓�n�$����=�ֻ�D�Y�!$��m�fO�=��|M���ʩQ(�*��N�9��k3V�`,/AV��6���@�d������x�y!�$����h��Aqbh�e:eK�����sI���.s�l���>���b��=���@�h�BI������Ԟ��=��BI��>]��7��:5�^{��|�w0Ȟf'Ϗ������ܝ���s�}�׮r!Ǥ�i��$�����+8L��'�>na����D��@��"�� 3D���",J'+	�V�U1)
�÷�{�U�����u���l&���@� 	 y�J�s8W-e���K�j` I����-������<�D���[S�UH{E0,�+8.
���H�
3J�`