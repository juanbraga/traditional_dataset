BZh91AY&SY�D�k 2߀Px����߰����P��a����ksp�hI�T�3S�~���4�OPF�A*i�<���F��2 h 	&��4����H�M!���M ѣ4��A�ɓ&F�L�LE%=j�h#�()�� ��Ey�"H-O��]�7�U�:�C]g��@W��m�CAV�|zO���Y+3�����E3������Iɿ����1w#ШaTD��-P�ʄ���[�ZJx���I��FX���s�6O}�θ�ci�
$v��<1�&�L����!ry���h�%��I��ibV@\�'�M�H\��Vc����e�-�FMrc���K������ccosm�j'��jy�p�R�d���VQ��w�ֻ��$/�Y�q&9�����t�10��&��8����B��ּ�w0�F8�~5m��Ϧs0v7�7�{�3\X<d{��׼��W盶!	��@�=���0]zġ����+(�я�;�ou!��@lP_�B��mz���D�r�/�Av�^hԻFi��=�c�3��ce"�f/�D�85�k�kpw���OY}��/%�6�U��",|����lz��H�*b��nj/F#Ft��E�yXSq�,?^Xc��Q�&T���e��w�� Pc
̋.U5m�M���07e����@[ȑp�O:��b�y��frs0cm�q����"�p��JV[B�g8� ��Z�r����AY�h��(�Rl$I�����JL��'	��؃"ȩk�b�
g�3��AP][�{�q-<�T�/c@�m�].��P΂��� �a^!|Fl8�cEc�V�-��pZ�Z,��UN�:%dF�{U�QV3��Y����C�1锪��S��:ä�!�X<�ї�ƫ/x8al�����R�2j$��(Z5Q���]G�H]�)�ؠ��:�®�̠�^1j�^�J�����C�QR�`���-�E�DJ* WDuߏ���)��%;X