BZh91AY&SYD�� G_�Px����߰����P��ZY�Z5��I2ɣSɡ4�i���Pd�=&�44yA��z���Tڇ�=@ �2  "4P�=L�i��#j4� h���0L@0	�h�h`ba$A	�hҏQ���A�� ���mL$@@���8�~N�Ǫ'c
l �2�~)�vP,�{G3)�A{Vmv�{����Z�c�s�v�/��Ǭh�F������h����2�*�����h!1Ga M)ͨBWc�) �GNA��9�/$��ci��8d6E�_�.�;9B[�#��V1�F�Rn`��vT
�R��R�����%\��T�*{)p{��*�����2����.$�Ao���4�d��}O�E�E��2_,E��ֻL�0p[Q����ؘK���YE���Q�Қ�PP�&\}K���^��m��q�4��������~�n�,E�	�Ѳ�SX�Sn/ĸh��8�8��e��uJ<g����NS�|�#��r�j�#v�G^fC3�@ءk�����ݤRSԢVY�(Z��(k�q�%���:C�lJب[\�\���C]�׫3p��Y����#��{j��a�"�˷�W�C��D(U��3��2F�`�.3ֱ	�s%A�'ѩ�5��Q��IHEz�0w��+!�8{Ӗ�%b|��Z����%~;��q15d\i1�i�2��N5/�z�N�s(gfa���:�,���Z�i�d-F'��<"���P��A�B��5�v�����7$��f�p�*�"N=з���F�y@�S�����! uu�b�ͪ�f����E��t�8߂Y�ߞh'
j�]����J�� q��m�
W��e��KRa�빀o�:�)��m�0W�MJ��l2�N>�5�0�"������^�[[��Ӡ�YڈV^R,�M�Yx�	L�+$Z�mL��$+HN�,�6YH���0rAc�Vh�tr&e�0���by�3���3�m��.�*��a����9�2�)㎟���)�%p��