BZh91AY&SY�9m� �_�Px����߰����P�p� MsFڑ�$H�<!=dɦ	�&�f�dh5<��Hڑ�<��P0��  i�!T�T=&����CM�  4��0&&�	�&L�&	���Q4����ѦCG�4 h4�X3��%�Q�D�$�`!��hD�D1����I��Ṕ�!r�ȋ
�V�~�r��lI7lB��B6Y1t7�}�Ӱ]hx](Y�;j�!��4�ҳB
��L�NEJM ��"�p�������d���4hjPG�%}i�ֺJ�XUj�X3>A��^��Ŕ" "g�?���A��w���z��$�-��V��L�/сxlP1$��^��=�%�*��1e���U�6;� 0��$
#Y�w���Q�-�������ԛ��֧�� ��f10�jUJũ�hM��p*�.^�.�¥��В���w׿Ri��n�NeN�p���6+E�����'���/.~��B�Q�t3�~�>k��jYd�E٨��H$RIN�]���=�v�ya-�o9-�����ƴ^�Y-e�@@�i��H{$s�ѳŒt����Ca@��=�@�����il+v��U�pBI���o"��$�[�TSeW9�M�C��f�!o_{�W�A���!n�i�m����2�5�U"�W�e�8�Idn���e�z�a�K�,c��p���p����t��RNQ4�v�k�u<Xy��N�N����"Y\��E����h�db(��s�^1���܍b���vd:��'k��:"J������Ev������8���!ڿǠ���߾Z`������p�d�j��t5P���%��i�����5�XZye�,m\�_��
�P��3LN��h���g4�4J�FX����^R}km�Z��~����'"�Yi^G�.߽0@� ]�\%0S�e�\8n����^��<�24��v�3�i�
�$f���8�(���%��TV�Ɇy��K�~�G�	�]Re@�!��9nW�`q����Hu
r��$��Z�*����)d�ĳ�����_��Y���[	�8B�#)@Υ2��M�܄ ���7�9⋲:��d.i�5�V8m(�mC0zՌ���0���B�� 6�A��ZhU�N��F�2y
��)FRңa��簎4B%Tv�_�w�[�W�!�1���@H���\``���MtEEH��
��U�4���=Y]�de[ň�c��4��}d�*��Lks�R̸��rܻ��id�2d�V�������)�q�m�