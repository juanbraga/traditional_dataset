BZh91AY&SY�Q�� �߀Px����߰����P~\� �ID$Sh!�
g�OS�Fi1�(��=T�       ��!=F�z�����  OP���&L�20�&�db``
�M I�=M��m�   Ѧ�`A�y Ƣ0$%�����W3�?��,)#��js�W�?w�4(��fG& �2Rb��ۿ�4� *!����2�h��E��`	�'vw��M��%#�2t�fL�ul'7�9E��Jb<T\ά�ʆd�&�������	F8� +��\��=��L $)��������V�Vj�M˅�q0���T��ɫv/&�����S�xL+�6D��[tBh�!Ig2��ω�D "\"�0'��Xm��2U����t|���2����U�Z�༽�Bt�5"��\�`�.�/�*�\�Bٱ�W4��C2��[�i����|��f!�`0�P I�P˴��h%�jQ�-���Vh|\d��Yy�fW��Y���a�� B���Z5�L��`��{m�����	JB�Z)�6����E #e�xO|��E	]���I		.$�"`��c�96Z�",�4H�ې�)N̒��Z2ږY]4Gʑ�HU&լ�N�eL�\����(�0�8 0���_��m>er��Z���1���{|�0?��Ň�s�ٻ��� �vϯ���@7O^ߟ�/ 4���<ݔ<s�l<��d���]Ir�=}ʼ�C2 >C�����std�ۋɆ����,]9�׿:�'���z�I��Ne�L68���Z�`w4�L�qk꫞-�zNW�N5��wh%��g�P<���2��L(�ص-u����O5���gm1���U��;A#�iK�7�ү1��A0�� ���z����(�6a�/�
�%�9�ro2��iL�\?���� 8�����V�&���8�����b /V��0�[U������u�+.uqӅ�
݀��w�6���\|r�K̎l,j^f��T�YZXb�腎Դ�m���9)��A3�=Ο���v�<IT��	����2�lH��i��W�xV��F�p�9OnK����Ő��ʹr�fԱv}8;�꣹5T���rk�&�
���*aVl;�K�t :�/��f�ݜ��q�1�eB�}��%U���k�E��ښ�Ш��S.,�F�7���K(ʸ�l��6I��yz&���.&����3��i��X�GTĽ-���+�KB�htP׋��b �2�jQ���?l�:�.�L��+����w$S�	
5O�