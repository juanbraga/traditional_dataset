BZh91AY&SY�>eb 3_�Px����߰����Pq��l��hI"h�h4hQ�h��2�Q�=OQ���LOP���&L�20�&�db``�!!=S�xL�M=&�z� ��0&&�	�&L�&	����CS)���O"mMz� $�SH4"BH-O�|�Y���d5�t��f
� �G3P�Q��6����p��:?C�%�YO
�b�#�{D���h&E»�v�\�\��s���H�J�39D01s��&���^�䨄�2~��q�R��,g���E��Xў�V1q�6�@ɚ�Ab��`%7(ɇ$�_G���V�hJ����}~�����r������@��#��cG��n�Bd��D�="8[e��%I��A|9A1ܚ`�N��Q4�L�P�Szإ�qw	d���<�d��[ o��TVr����v��NGɟn�M��Hq�GO����T�����v8ǒ�!4�,�S����Q�;�cO:�[�m0�H���Ǚb��u���*`r�\�7Q4�i���ŉ<�.ќ]��Z<L�ro�7h� 	��~���e���W�#}*Y��m��̖�3n��aӱ�%��FE���)q	;�VD�4)�F¦�#���T,�Ԩ1��2�h {��+;�6���;������00��*G�	����P��Da�D�t��Ŵ���NAa�@�b�Ɯ3QT+���fp�*I����Y����D砱�p�� �-��9E�%�ӏd��^<u�Z�2Al���ĕ�&$��B�Ĵ	 d��$쎷gZf�V�Y4�e g"�	�y���56}z�l���R�M�bπ�'��k`�d�8y�oΠU�O>����N3=�1[6p�e�KZa�娨-�9l�
M�JE��2P��R**JhEFq�a���r$α��&xº��~{/=䂾	��%f����%a�a6:����1F,��0(��k��]}w�n橍E�؂f�@�Y��)���-�u�֯*܋啹j�^f\��s�scA���^n�����"�(HU�2� 