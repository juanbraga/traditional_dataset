BZh91AY&SY�r� ��_�py����߰����`�>�9� %�(��Q@S�         !���T�x (�    4��� 
d5��#m"i����.F�[�֑��wQV���2�9ΣЕ�F�iP F +Fk� H2b�R��F�J�����Z,lT	44�  J�ذ�(���a��P.��j�Ѭ6
l���TKa�0 4�%DF��@)cT�%*$��5�"�l*I(Q` ��cJ��T�)F-%%J!i���iF��+%3�  X. � �����@P 4� *�Ȓ���a��L	�0 &2d�L&F@��M#4i���T*! b4d`� 4 114J  �������=&�S4ɤi �*�22i���4Lj0�_=��]�+ÍkKS�%�q��Z(��"��UJ
�+�O�"��D�>����"FH }�Y�g���U���@�	&�'�BT$G��\"��
�����f�?��0��aT!�RH �2 T,���B��A@��&0�@	VE�!R$$X ,�R@��Ld �@&� ���HAH�
�* � *��$b g���C���C�'ޝ !\DQ��}C>_�����3�%�&c��j�#���N�CIv���b�-N`TLS�*HBr��F�����g<�h�jls�y��\����uu1�Wy|�����	X��3u�� �4՛E�[��R���T�n%��^��K�n�HٻY -J���6��m5Y:�m�1S̏*G�k4�ʰ�l-�ti�1j�X��Zn��n��j��n��a-����0Q��*���[��f)����R�a��Sv��~��2����&i2�2Mc2�,�0��vN��y�]:DA���öv��)�I[r�0L*D�VjYy7X8�ݢn�U��i	���Zōy3�4�«U[�R�h٭��j"��vЖA�{�앗l�QD��t��*����v��D��V�ToE-��T�<�d��ޒ�'�jm� �x6ޔt�b�mf�f[�Z�e尅�؉+ю�
��Q{c�J
�3R�����k#9q.2��Lw(�4 �Z�1��q�0��/*m�Cjiմ�'���E���5���Xf�^&r�>(Y2�THH�(�Ç2j��W�Sq[W���^m+�8=��f9�spߔ{��dXa8�x�x����b��QEb/-Q�E��)��UX�AT;h*�X��o��Ǻ��GV�+R��.���ƭ�mQv� !���R���i�p��[��JD��ni�G%k�u�̽,����%]�l���/
�L3u� � �OJ�FTKM*ɇZ�!�6[�T���w��R��R�l��יe	�a�y�E�2��89.寪m�'�$�QDZ�Vt<����Cs�o��˳3�6pE�tJ��RX�җ�+fƕ�E+%Z"ÕbhŶQb�+K�z6ݸN"��0]<��8X$�1���,���f�r�U�����d�%B8p������B^,�N�G+kDǃVeú�h<�90x3E���K����J����S�ke��W�����t������#
yW`���qYq^MZ��ô���0���5hMut�f�e��0/t-<��������ճGc�fň�4R�wX�3�[4�����di����e�Y��)�)t�y��n�b��!0������a:�#��DD5�'�f(m�(B��0��(4���5]<Zä�/ڝ�i�$J�x�(�92��}�[-a�A��۲Ac]�A Z�Z���l���їRZ 
$J�L�)<����� 0����W|���G�K��--%y�tt�o2�$r�����	�!�4��#p�n�5�LXj��VE��U!f�Y�x��l�j� �`�Ð�I�YN�:�͚�\Hl�J
R�V�*�
:MRv�w�Y�5nd�8��HD�ذ쫔�ԝ����U��b ��XNM�x���IZ͏,�S� �A+q2���*BP2E?dG5M{�!)�J��F��f
d�6�
C;Æ�����ުt�9���*�Z��v��5�Z�R�A��HBT�3�q�(�hWe�I�P���H�m$DW-UM5����"��z���j�A�[d�#�	�yi�NʇF��Yp���^�y2��22T�l[R`�w��67\��Xb�U��f�j4U���²�,9�&5���gM40]ҽ���<���
)V!v%r��V���K�;k�>a]��0kӪؘ6羌%>����5���H�n�K�+HZ��������k)3p�	�h�^V�M��ڀ(�l�dv�X�6�
�ʹl�M�P&��V5��\����Dy������͸CBV�0����r�\�Q0���9��9vu4ta��ͬ�,�Aл��Il!�*]�"���ʦ�I�Ķ��41\PN34��o-qo
���]u��ki�#i5	���73.�`�u��(�Q�d[s�p�u�sS,��0�h�(Lh�˃�C]N0�0k&cR�i�-m����XL�e�^"��弥\dsih���z���Ժ�f	34�M�U��-эt�D��[,�[��3qsXRc�Z�46bF HY�Ui��.�T�X�C��lKH�t�l��Қ��5�R���\��ҙ��[�
\9v`�"Ei@���v4Ɍ�f�p�f+����ekIx�m���8Z�st��h�	Ħ[�,��6εK��ڕ50nb� 4V��`�G]vWE��)[u��b��5t,�q.�
��붚�7U36�kI`�ԍ�G3\��M͊���%�L.���<P��Ǒ�ر�h��%f�b��*T&�4��� ��n`��`e�\gL���i��떁n�9�62R��R�0ہS:�Q��%IM4ȋ��ЧkX�Gb5��k-���\����pC�±H%����ZECl�lc3,����7KK�JWl]���噙��#Bm)6��G��[[�f&�6v��0�J6�� �m�%.�3
�5t�*�7D��їi��l(د�Q��#�l6ƈ�R��nie���+abX��%��5-͖��iYSr�s����7.�8�Q�i�A��sH�	��\�8�jm5�myT���-�qWY]x�L[F��2h�@�M-%�o۬�hu*��q`�l!�}j�:�
�j�$���(՚�s���ny�fK����Vn;h�Z��0�W�y�ey��M)��Ժ��	.
UY��˦�4qJF&.�ʵ��1,�[��`,v6��&���Zҗ�KE�f�b���m�;\kf�����uI]en�)l���YNm���ܢ�-e���6t��FU�F�����+kxcl�e��`;��Z�\6��c��B�AȺ�E�7��GnjY�-�ĺ�[�\��e�ї�x��%����L&ej�m�������ٕfSK)ko���6��Pa]�Ԍ��vVF��Xe�eCL����d��v����6�\l���B;f� 9��1����<�qͭq3���u��5��R�t5uJ�[Q���	B���k.-�]�[+-j���8p�r� �+�6��M�@Eq�_���{i��{Yi��MG�+� �<C�]��S(�;�&���� 	I�R���9D�"^*��@+!�I2O�I6�<H,4���$*B�`���`!ԒI1$i��d	�Lx��&2��{��i�U����6�a�y���8�!����=L���^@�V�P1\���:Q� �!c2T,;?��d��V�˩��[���Y���/C2�������'�W�"S2g,%�R���a�����jqJ��Z�V+�y-T}ǆ��C˖*ɔdK3.&L���[�f`9,����x�c��ɶ��շ�Z��ASf�b�1���d(Tif��@۶uU��\F��e�̼�E�Kʳ#/.�g]����T�5�Q�\��C���@AY!	#8x��:�O��O湊e����g�9RS�e��"��h9�--
�N��L�n%l��([n��̶a��D��,U��
mn��sV�fQul�)�s`��M6�Lى�ٝi8�\�B�댶��lZ�B˥JM\��F�]��BWYm�6q�Xճi�xij����%�A
̸%�-���i.3fƠ�naM-�YAn-��64#o�"֤n.3�\V ���M��D��'-��6�Ic�����fR96��$-�qQ.���N)i��LfŨ�-��ˑ�������n��Y�Qʺ�u��$���!rN��־Mw�Ή�\�4�T����j��5b�MV�m�f�J����V�*�f,�ܚ�.�G.J�s\�y��@�H����".�P uD�@���6���C;B�eU%V#ְUDX�DP�ETb�`�
����
�� ����
�ՠ��E@Y4�	�UdQAV�A����EX�E���-EAQD`����u�U*DET���A�.�UR(�E(��H�TUDAE���#��PU\޷͜EE"��0U��PUAV"�آ�+w�
�b�Q`"����R*
"+�v�F1GV��*�����]�1n�Ub��T��Fq�EY����E"��[�L���X�zՌU����^e9)EUE|j��b,F��Y�(�z�b*tB�J�X �db#Y,DTF9��vԘ��V1��T��mE�����4EQ�2�U�h����AUTF9j/�Y�(�EF"���Qb�����^pX�� �,U���F(��"")�QdQDQ�
�M2�X��Z1�U�U��m낪"��n�X�*��Q�<��6�TAA\nYF(�YYQ"���wMآ1Q�(�l����֪"
�#��Q�6�{n�DTb�ETU;��G��4ł1��Uc-N�z�G)UU���w}���hU�f�ݗA"�yy�z�>�As�`�"���X��UL�~���L���<�#UX���U��"��>�|�
bT����Us/��1E�=�W`fPUAF=��X�ח==�y�~ִ�
x��m�9p�_�?�$$O��2����E�Ԫȥij�,Tc�E��ZQ7��)����洧YE����_|f�(��.5E�FбW�Y0`x�E�YX�h��n�<͌XǟPď�U�,Xow�W�i����E�����A�Z�DUP�Z؞�0QF�1�EE�*.�Hb��W�2��J�(����xq���`�﷚֠�LX�fQ��5��׎�X8ب�}�s�����PG-g�Lj_�*���=�{5�c���K�V����_v����H��M�"�{���2���y����;�tYTeCI��)Q�t����'��"����8*+=J��d��z�DNeÖ���A���c�.'�\t����ѳkE�*Kۊ*8�V ڤ �RÊ��b����QIA�4�·|ד�c30���˙�b*������vu�D�֨�p�-~�x�G����3w;kݮ����ØV*��廰�W��Ķ��~��V ������3*(�.oKK;�օ�m
ֶ�v��3�̱E�"%<��_.:[�n�]Z�5�-��fp�(VVhCߵ��1��i�Y�h÷0�����mh��q�*o�fj�^[�����:�Q;h�r¾�otdSi_-1R��Y�YKue�ˉ�S�xq�E��\�c^�4�����V
�0=o)�Wm��yq�Ugm��V�O|��b!�1�̾��_n}���X��ψ>𨩓�pW)��:���nk�DS�U�߯�{�$^���|�A���^����^5�i�y�[�0�%���[u���Ɇ-V�71r���k�e��g>��#��Z���F��������aآ�w��>�������kS�Z/��T��y��~���u��c/y��:ɾ�B��k�u�
*��b̦�~tbC��G�F�	��
oX����<���I�#�`��_tΤ�L޵E
 ����Y�<�#	q�7�죦�YG�փ�S���̸()�~�9��--�`^�Q~fןz��N��M��M�Իf��u3e�630Lk.���K4���̫��űv��Y��a1�K`IKNY��#@�	oSU֮}���� �S7qF�̭s���Ll��~{���z�\r��nJ�l�X��v\��D+���e������s�
>]<��>s}�V��Y+8��aĮ5y��oP��ܫ�~F].� �����CZ�I�EaS@Q��&
��-� �=�쉀���毄:"�`�M������߉[(��ɰ��[yie��^��Ƕ��9��Z�{��2q�-�S�p��%�d���Ԥ�>q�>��r�,�I ���3�?i����iq�^X&ز���w��`�a%ş�7q���,�
 �1 
fEg��iU�db܉���P�܈#�6�&�
6N꺤��7ۙF6.����56��ۆ�S����MD�P�
���6��}��w�]/Auf�9ЮZ$�9����ƿ&9aX��{��U�:��u��k1
�}��g�5�3sy�yM+�1Q�bB�kd*)�b`" tu#H����;F~����b�������d�0\�Uir�
y�L����nٖ����0ej�x��8�3*>	�H@.c�-Q
˽���(��7&̘���<�?I��k&*煮?}���F�}y��+�M�9@�r\��{�r|��fA=�+(�L?����V�ᯇv͸HΤ	F�
��BM��e�Π�ʼd39���z Y�$����,��ZP9�Th�e
���#%�a�h�*��a"��fF�c�|͜&�c!��庉�`ۺ�S�jX1,fDV�4ځ
�r\`��Vx|+���4h<�϶y=����wR`ms���^S�/y�ݤ�}��Q���`b�L�Z��b���d?#:���0�)�]B~����!�
���Av��Ĩ�g�"Hd�$u=c.��p.�4�ӑ�L�O�x�p��ekbLĿ�y��Q��"��;�r���U�f�7X/b�JQb`�)Ĳʆ؁
 ����M��[H�,Į�[-�$�Y�eb�ѶhW���R���Ţ�x�h��S��K��4������dD?fB�A@Pǲ��H������8����uG��U��_��^W�ӝ�+���F�G%���'�)!��*C���|�rF#t6\��+��$��:��
##%� �m�I#�&��Vc����y�2��c%E�{}�[u��� �$�"+ Yd"#.8��2�L?��u`�\U<��e^ְ-�&�c��H��L �J	���5�T�Y��*FS��5�dhၤ���R1G�NB��P�3��)4,�"�		�"鐁����.�|0]W3RWe�����z�u׶o~��<me�R��1��~2MDB%/��Y�Y�I:N�ɡ���2Q�Rj1Ԕ�a�!#��q� nq�Q ���1n6Ug'H�?C�~�S���Ʈ��1&�R�v&-'�""0����pG7�S��M�}�\���Powb9D�'H�%A���]+gm�.�8�gNP)�@n0�Gu�����A�;�.��Vs��i^^���M(�!.:i$�t�eѰ^ň���M�ѭ{��lc-��A�Z0j�����mQ�[�O2�8㠄Dx+��5�|����?-}��x�&������ȲI'��b��"	���:��Q|�� �D���=�	ր�t��Õ"�Hb�GJ`��DG���(Hq(YkU6m}�g��t�{R����Y��\T�k��4l_Dz��I$����I�Y3o�(�m�,�f/��GJ�WԨ��?/��~4Q��J������ �n�tap�DY@�DTB(��G����M��i�y��u��֪-~pG�Ly�j?������
��Z�~�m�E�Q�����Ug7�)����S��U��$�D�[�(�D�����tB>r/Z���ڣ�O��Q"P�L��3�qN��$�u#7�h��|G����T�7�Hk�LQݮ��?�Ŏ�E�YBf��e|���o?7�v�-YGN��Jc߱���iV'��#��)aតD���	�=;L��7���Z���r��7�!�;�x�K�j~��	2~�$A �@,B�}��ȝ�b��"�"[�SL��l��64��$t̎iZF��'K?f\
(�:��t��?A�	&L4�$ؔa>�S&��aD�0�B�y��q�HӀ��Ҿ�C�
1� ���T  2A?+�}���'ǖ���l�,nǗ+aؐ����fՑ`R�WI e5��v�I�Ląѡ�`�R 9�kf��hK�01��`K�a���L��&Yc�ֵ�>PD\��z�9Co��6��NJ3�%�@C�|�>$�JA�N#d�T�����=��8����y���Y���3k.�T�=���`>�� �<}h#F���1������y ���yJ΄��ã��e/��l����ݻf;���7��q��wJu=q���8�d�0�O��j��B̞;&�~Kiw��5=|ʡ�4m�nS-�i}�����ϟ��O��Zmr��c�5�)�/�,*e�~f�\wW�o�̋ޕz��9�>��<�S�^�UE_��ǳ��3"FJ���w�~X�>��4��+_Z����U;.�;��R4B?"���@���F���������]��w���u�����$2 ��@�_�BC�����$
 �+H��[xdmG�ÛR�<�,� H�KP��f�N�v��6J�D��-��o7��!�1�"fHl��1/iI:�l�r��1�q"�|��6��4�`��B!�r��B���X��tn4RD��g��R$a�e�'�fy�����M
A_
"��R�)�h�p��0@���#H�u"H!�4��4���W�O ��%\`��V_�������TI ��B�S���R��R$����
�x��^`�܅Aڈu�X"�Oo,�m��H�m�2E"jc�.���FOȒA ��	��a�p���0���I�/1H(��i^�O�mU���R��Kj'���vk��f\U|aN4�e.SZ��Bha��<q(h~�؉�z�+��[�^�UWƸ�k+]8���ǞX`�\�UۢB�3���Y�^Ѐ>1K���_Y�Kw|ɪ? o��@����&J&I������@�D�Pd�z}������Su\&F\�I�t,��87B��jJ�,��|��blV����n�|�|�=�2�V{hV��fi[�N�K�6�J��c��?r���	
��@�|p~�U�
 ��4�����{h-o�N���bO����� +���/�|�-54Ǯ�qP��	V�Q�7�$�/�RQr��x��(Y�~r���
Yzb��;�R��u1y�M�ձC"��7���%��RV�)F�5�I��4��0��-��A��u(��2.}<��|e:>��y;�[��ߠPz�|=�5��q}��	>�?�MM�1,�ߎ �H��0!�o�M-������j�Y�̬��@27V�e|#��uU��w�2.�k
t<�Uua�\��o#k�/��P��`�5@a�Qm�3�I������y��ex̄c��J�Ҋ�K���ƞ�F0t����f�̤W��*�RNJ�%Ұ�U�X�PX�4���X������vЎ��f��@0;�w\O��0��}{��_z���l�غa�LCHxB�Y=�*P�_�-�wُu�^u'���S:��X� ]��N�}{u��T�{�q���G�{Z��Oxs"�HG9�F,Rzq#z��f�d�2�:@�b)?��f>�͈;Ľ0Rt�ߧ��d�黐'��Iy�;��Aj]nh�͜���}�H���F)ۜ��/��{fH�#��b�$w���[�����eo5�S�f�ɉ>�CH�[n6Cٝ"G-ˀ0�{q�ά��q�5r(F��3&V���~o^LQZ��sq����ל��V9�G���b��$WM9�ywa��g����04�66G\53ђ&FG����Rǜzs�/�K�@ˉ N%F�3ә�����h����F
�8��ZU��$��>q��A,ňy2ߞ�O�ݸ�#Pw����C�M��ĥ,d\�STT�"��ợ���C����h�\��;J�D���;�Gn���0��L#�:/C�]��1>ݝ�:���*1��+z/�>�m�<\ �p�v�9@����MiP�Y%rl�|ԭ�N��
Y�k0�w��CG�H�gN�AZ�/D���6�7FA��<l���E�����.� [d��*+é�ق�[N��}�M��Z���sMn�u���o����kT6g��.���18�dC|�$C#nmnJ�6��4� )�I�[��q����n���M�-��[�K��������v�X�!��h7e�ԩka+�JmR���QɯъJBjՎ�`"�Qf@��ـřA.��f�J�[ۊ]:UV�]�*u�Ԕx8J���(Q���,�i�J��bK���v̪YZ�d��3�^r�.\����6h�!]FX겑��b��.��r5���G�nF�iV��X��l�FM�����gg�	zmxw���1Z��t�Gl:��1���lr�E*�ܔ����#�c�$3� F	���K�9.fF�l��_����\`!6g�fhbr|Nn#��jq�1
1?eɝ}3�3��Z�Qb��$�.EvdW�n�}�x�d_����YL�z�����ўD�s	q�Q�;�@��АE5�/^P�dl4b6Qe���%��O�vl�G�=���T��̦4fP�	BׅLF�U��8��B�_P�I&�m�Z#�A#��)�N����+҆�v��1w�J��S��m�s���r\q�Q��˸�Ϡ���Qq*��#�VFG�����C]?���]�r�
���8a��a��
ʯ9][�/LZ��ў<}�6�	�O�oZ1��^�le��=�r���*�Ǎz�ۑs;�����e��2a�&�i�ߊ�����X�W����
���(D^c���3��`���\}��m�y=��OX�@�\�r��@�C��;]\�bWޱ>�d�>����.!o�`�8�(�X6/���^O��5�'��1=3���� ��b�_5n;B����_�m�Z��y=�#�^M��ax\����̂�Ry�A�_|���;��ZS�٪5h�l�B���C۳D��R��C^A��Z7��0P��\�r:��t��ꢭ}��QG�y�&��@s|1E���k�jSA'a�ɏlD�k}�e��%�H��ʍ���B&��)�_1}a�޻���:������0jvV��͕Q�F�B�an���W&��A��i�W^kK��;9�4�6�h��a�6tU�_�C�!��-�!$E1�w�Zw�%Ѷ}2,�6��?���S�>N�yH�N���-Vw��I�?�~����S�}
8z#J�wXv��Udw}��k.�3�ʾ�8s7~�{iǽ�1/�����=<E��T&8��-�e=왚Pߘ��ȚW�\��
��9�V�D�lov���cfƨ�U����vPU��G� ����	��c�"�nU�K
H蘎7��&v��XI|��+;bC��:�+1�A�HU&��M�^i�����>�p��-�	1.J�+�d�I�]L\�td��ჲ�QNVby'*�Ǘ���F,�>>�*Ͷj��<K�hg.ݎ%J���#/4��-[�U6�ޟ�/b��U���
{3�q�>6�@�=�(\�ģ��x3�����	���w�����l0�pن�
�����f���5u/��A�>��wϣI"�i���EP����"��5f!���0�(T���Ж���S�2D�0�9!5'�hƇnY�ԗ]��祌�s�̨�dX�h��q4������@>fh-����N�>o:���1���q� ���Rl>6��"���02�z�5�~r�9P�ݫ�� -c&���<3=#N�U���s:|n�91ƒ�����G<�~C���xh'��]��ߕJ�T��yw�=_?6G�/+�)����Swb4"�_�4J��4�2\�u�R�	f�iM]��jhL�nŖ"�q)s�Y�c�ͳ��W���ʅ+
��H݅��f��Wᣳ��7�{��X�.�C�����!kMx�ї�0r�gf7�����Dw���]����0�Y|����Y'�'O��o����n�~�%�	i!Rf��\����XI��M�̐*�7�7}�r{m�ک��0)n�1���T7��1��ۧA�I�S���{}?RߗB P��u����ʢ�����#R�zqF?`�
�R����n�Z�!�>;�s�T���4q�}�Qdx��ۻ�
�c�M�J?%|L�)��_���ձq�±�W�s�}�LxD��u�Z��k+�������t_�/���hA��N�q�.�co��f��hFi���t^ܾ�4m����@l�B]��oG앹YR�ɪ��M���ͣ��6��3U�71�q!�	W/'q��	z��۝�����\�̺��a�7z�㦙Q��*Z0���e�λ�����w�,�z�ݩۚ�R�Q�kE����qp�Im<ܒ����m��d���un9��2�c�|,�X�v��Q2�6��кN�����*��hu/��p��|<�����Wv��Q�y�F��*tYt5�3m"�0a�D4x|��/﬿�:π{toG�ә����gK��_�P\�S& �I��/�-�.AV������#��Z����
���n�@T*�2Ό�3�Y�TY�Q>�M�( �PKm�l�Nc�5��Ys��9zd�0��8�q<"���z(JI!mA,��N+����NJ5�NX�@���L7V�cif��'0���6�=ѓ*kvD��<vU�*�^sOb�0��Ԉ���!,�`��
�Զ�, ���6f�̠��m��1���v�����͆ٙFVbj;��GZ�8I��m�c��a���~��$�����xM��.�*�)�m�y-ߋC���x���\(Fh�^#���|K�R���?&���An�W�>ט<9|���]}p*��X5(a	V�0b%�A�,"k�AZPA&b�v�\����Bgd{7�z�U�hn���@1is���O9���활.�pu[�nⱑ{�4�M��ㇷ{��w�Ss۰b��h��Q,�����
<9W�F8�Y2��F�����3|8�E��t��4mZ
Ց��aQ��g�Z�zC�H:�k�����w��#JS�{rX�ẍ�ɟTࢳ��ǯ6����w���*7�vo>j��q�]K�ȸ�=��9�!�5I�ɑ�j�oΦ;�׾������N1�j��|�:;�9�N�W.qx��f#v#)��g���#9�Ѫ�G<������=I�ﭼƤ������{�؝�l�R�!:��I^wgj�s�:�-E��7�a��B.V�>{a�Uy�T�Ezi*���s�}��З��>�ź0�3U�	]~�N8�M|0��&�
A��=8��/b:��j~L�����+��+�To��2���tT)퉢8ߏ(�JGm�0eŜ���Q��0�G���m��u�3eW��=�yu:K�a�ºV�P��q� h�N��$�!Y�hZ�h�h�驁���\���kij��T�2��n�gs&�g[Z�	�G6�mu*6W{ ������x�H��p���ҧٗ�&��}�&&�Y� U�Zci�f%��c������)�Io��ۻ�h��_ֺ|����i����s�=Fg�qO�5a�T@M��d����v��Q�]�a�-�J��t<]K��&�U�6�`j%�j���P;�j{Gz��DdǶ�G���2k#��Wm���.S�Ʈ}
�R�z��F@����D�Tݻh'*>�)]o��.S�`��a�ᶌF]X��1��L\�@޺3���,=:5�'iA)�=�� ���X��ًr�qw�3�CP��Hr��`�}v�R��օ��u=�H<�y
Miod"��ة�Y�{2�q���H��m*�{2��JvA�^8D}����FķuG��}����6|��v�eGey�����.LÕr��n;�ᰖS�ǽ\��͉���P���VT�>�K {ʧ'��}ǻ����F~UÝ�m"'�Ë�A���;}�q/�_#I�Qn;tUw@P�p���C�<��q,���g���v� ���>�x�&�����T��^������(-M��*�Ha�w����+���|��T�����[o�D�t�>�1=��w~3�ڛL��Ԙ�jR@P�h�ZSX_V����E�|;�?��
I|���sS����R�g��[�ve�Y����^��^3f�T���ɜ�3�Mr�ۘ]�k�==�t�v�7�spL:��C7]��H���*n՘�TF��[>�\�7�᜶�y��T�����؊�H���.�3���s[{KT���;��s�{��2��4	{�)���[�5,��k���׆(�iu�k���L�Wf�vp.L1�׆�)��-�-��qm�^��ypj��˘��:�	5Ź3�Sl�i�M[R��#.�f����4+.����p�Fm�"�!�W]W�Mo-5�.�3npjLD�˪cf��l�Cl]��f6��K* ��nfMy�]��[Z�5�-#ln����Z�G]ste�XiJ�n�e4y�m�n���qYq4&���2�����'Y	n�9������p.¨XIe�V7�.ZMt����ӓ���N�W�_,k��K��jp�jkJ�8�[-�p�̖k�u+��b�pi�kei]��E��)��j�����X��T	��s^S���g�Qw�,�o{j�^?������T^��v��u�Wc�Of�Ļ�g9l�5
��D�f�>��IN\
[Gse�<����WJ�<��ئ�k���;1լϫ�Γ+�l4�p�p��� ��06kgk/������QR�(EQ��VyV��]���P���,U+J��F ƅ�e�xk፭l��5>��g~�pO8!�46Sq�T��5�Z�w��B`��b����"|��h�T���*�*��ʒV���N��Ϭ��h̵��i���K>f��|���#�һ[���_gwz���}q:@A#�K������4��B�(����J�1Tс�d�/?W��{V5��T��ӌ�-&)���M�h�jM+����;^E�A�V���dzפ�ĜY������}�j���;�ǐ��o���{P9�y�pmQQ��]��\��v�s-�IǗu�/'��ߒ�o�O�&��l�]�gD�ޖ?{�g�^���a��ݛ���F����#2���͙.&��Q7g��6���v}AQ2�>�.��T��GN�#�ɼ"�F�j�8��6��&�~q}:ȸ
26�y�V�@ �V}��8�"+;�*��jB�'�<�����/��A7�SL:[�eq]��q"�b(憲�eT���+Z�r8Ѱ++Ű�]t��-��M^�Ҕ�.�Fh���3wڛ[I�N{X�a�t�\;��M�v�{�^D;�L��(����t}T��k�b��pe�[���p-K�2UB�𤋮;^fOј×o�{��{�Bw܊�w�.$� aÃ�j��3-��{'�eg2�>�*^ན��l�	��1]R��m���*��)����btF�[c��[���y"�^n����~��RVl1P�b+�
�q;ݦAD'�����U��R��s��6�~��py"<87
D(e(l��1��_M[ċÛ���)�W��l���>V�]��{1"����7�:�SU�*Q �#�no)%7Ԣ\;w��0L��P����*VoH]�vj��w�eҊ���T��;�˨F"%G�=ՠ�T$A,�B��(Cq�?9wdN]��A��f�"��Q\5]EӔ?xC�+v�����W,���꒣��v'��Q�~@���;>Ж$���0�ӹ������S�>�AzԎ�+<}������8v#*�q���m2�� �h
�F�%J��Թ|���f`�G��'ؔù0V��q��:�ݞ"�mƋ]"�=Hf�N�϶m������Z��۾��[�������e!�]}�T�N��kߍ���:�p��+�E�o��@խPF�m��8������\���n��	)s4�R%Л��Z��s����Z�ٚR�jIT�يk�J&I.[�O5��:�oκ�'0U�%��gv:V�*Z��|2�f�6pQ�Q���@�\M{nv74z����M�>2x�[�J�ߍg5���`G,Z����n_q��1�X�a�+NW<ɲ5���ԞSm����if
��k#G��k����c(S[��9�hS�sB�w�`��f��"3/�Κ]~��ؼ�	:bxKO'm�;�I[�}��p����d�\s/�{Ev�]�}V^���>q��E���*�4�V�m�0Sb�V�3#dN6�xySwT�6/�\h�<j�t˘}.�⯝�7"�1T���/FuO ��V�l��r�35��u3�63�c�o��q$+����i=W�/��P49��T��
��+�	sW�|������a�4�)ё��������(�D%����#�3;H�u�K�u�u�VJ���I@#�DH-�زF5�/C����U:��h�ĺwY�Nmq����Z�?MUS4�)���ǸF��#Mғ�W�&�����2��Tۏ�����y��l6�4��c�����{凩�:�&�r�����Ӎ}��n��OY�0��d�m������u˽�{���7��k�R��>�z�r�nD���sg�{d�F�6�)����+Ov�e,`q�K�RZ��vެ;�������r)]B�!6Zk���A"�̴���傖ɗ���>�����vn7<9k�)G91*�l�8�����ڜ����Ҕ)�u�g�tM�C�~�Rd�ʃ��k�FN��6�b�Hm�.�˪��>�N�>���O���y�9�	�Y𺬳��	f��������n�<�̈�U"��������Y�U���~��_&<�Y�DK������׷s=q�@�͌��@!�qyA�ߩ]�?H*݉p��y�^�)��o�u-���l�Y���r���v�M��fք�Nl���V4�\+R\7����4��kt��)�M�l�l�.pPn`\�KF����f�,����df*�U�;�����ߛ�{|��`����Eׅ�J���g��y��2~�6l���
��U`��q��&Ek�T;�މ+9�pę���O��qJ=3lg	��DY��W8��r���|�s4 gi&���h�����}��Y��S��9nl¬Şq�B���Xxs4���3[������ɭ�~��hP/�	���eĠ{$Q��������h�'�+��4Ky5�[�� v%�o�����C�u7S����CMX��!rP�#���k4Rˬ�Ό1�����hD#����e|���y!�v��o�QU!^b����b��	M�Z��ҍ����;5/
�h�-%����K�{�}} Ǽź��Z��n�lD!��Ap�JP�!�]Е���vk�7J�$J�-k�=�#�~���S1#�o�����s���Ӷ5<��t}���Ƿ�=0����ƴ/N��+��3�d�uVm
e����fLb
p$9Fn�<��3��W�)�۹�Y���(m4�D8I��m��n��B�<nH)�\;.��XJ�*=���`̯f����D���L��=��Q�A��L�|���l��}��6ᔵ���b�EİTԍ��qF��}�u4���傦�<��	��5y<�t�򹹙.�$�u�hm��n�s��M].�B�����Ɔ��]��R2b֗B�3x�,.�c���10����χ�Sȫ�.Y7]��h�v�f�vn��n%1Bӝ}��0^(ЄT��<b��x⮕�I���֑#>�m,ށ,^yX�l��K|�Qg�G�����N��	�	F'a���C�ۺ:};���{�.#=4`�R��M�.g2����n�9�u����S� ���V�=z�.��q��h���B�ܲ=�7\�8O��|8zj��>�Ѫ3�s�~�I٫vм:��y��h#L���D@i��GmKT�7=l��ً�A�B��j����}��R�K�9\����v��a"ēU@�ЍT�.!���<Iu�-<Uz�_��z�upE1>С2���{Ǎ�Hs"�/䉇�L�h��w�2r��{0��|�l�o��C����kq_D���B��~d�'�C�8�\~��н�e�|��R:ڿy+E`�XKyH�z[�ќ�����,��n�ں�FB��v�7��짛\�ʰPр��~u<|iz/���u��+C��`ޕ�k0h�,�3�a�� �{���l��)����Dw����U�=��7�"�l��b��%�ZA��y�b�$�S���W�,L��khx�0b5P֓�ULw����s�E�����ٳ��O�O\D����۠�&�����l~u��+gj�R,���S��1i��)A؞�O���߫�ᷦf�ˣz78���� �cPxlJgiŃl%{Y���"��s{r��J~�:�k��&d�w���z-딅)yJ�t��_k�I7���Ѥ���N3� ٶ�h�Ȗ5�����ҕ3����Il9k���5Σ��5��,���]i�b�W���f�V�r���%�k��pxpi��Ֆ���g�Vʘ�ic��.K� ��EIh�h��5d�Z���6�j��K+^�S�jm)c\���0�svԘcqR\kKv�a�'3l����ΰ�K6�Y��(��XX�K�s�	�8:��mK*��ddB`m�a��^T��06�0��f�m��J0��+�+�]F�Vm�7)Gm]�K�ݜmkM��c�5�kK�$��tq�$���<���`!��EXU�,�2����`C�9��ܳL�5m�)\���3m��&ZE�F>q
D��Z��o� ��TV�d����&N����=;$V:�s��	���cOL�/þunZ��mΦxx�����м�F<��`�f��1����ۆ�-��B(0�ޛ��K����#��P��u�'��d���I���Ⱦ�͡ik�=ﶫ=aƂz�!ܽʗ~��Ⱥ�����Զ����_w��;w74��k�Y��als�s璳1��q4��~(��	�NЙ���&g�蹬����.����E����tX<���;=Y�G�w������u��<�g�%�c 1�EZ�R�-Qz�s;�٬�g���P ]q�W� +�@ZFͤ�IV�]��Oi<�ʾ�������
�g�2��8A�2l�r��+�[a)�8f�sZ�g���r[�m�b=��;b�&5�NtJl�C�b5����9�7q�Y2�O�/��U�n��
��I+����P�:��E���{�s��G�>s���C��}����7��3�1�{�Ы�{څI;7��%�,i����	b��wL���(��gb(J�ò=M��UR7� *����u�a����[�5�t�mn��Y@����ռ�h<Mc@�R���F]���@����ZKiG6��u~�|����Ή��y�G��}9��f��fJ�%q��\��VcXL�T��!��p�ś�*��KFj*zE��v6{�-��n��{:�m洗5�PDq�w��&��Ju��rk�s��G7{Ų|�'���{-۳�s#!��DRx��nS��>�+4vZ�z�FY��}͞��)��{<"60w;q�r�F�ݦ2&��Ź��gie&�P����ׇ�:��/h�D�
�"Ce�b�4F\�Z<:ϳ �9w1�cأ�n^�e.c�Ze�s�n����|b�׉Ǘre�7���d8�=�ٚ���m�d箫�4���ޑ�K���V,$���C�,#Aa�S;x|�efE��y�~�7"�����E�[�����oȒ|��my����`8��{��	�S�'Q�P��,�g�E[�ך��.>k��4�#��ƾCءZIÆ�
m�s��j�W���V�;՞h{ۄg���ۼ��Z�k�ow&�a~��R���L�F�U�� �_���1Q�V�;a��'���h	�~�T��2�
�E��<���cy��@��������T�Ŏ�-)�V[fSe`\�[x�f	T�T�Ze#�
]�q:~�m>4NR��'�kё��q�m���lߺ�����p*�bcS`��H����W��Y���Ȍ%�xJ��<��o�"�*�FuoS�H�uj�YT���j�a�8�Y�	L�Пh\vsN`3��]�k�����NL�,�:7dZ���9���nX/��v}}��(0fm��Zj�C�s���y���*�����f����,����u؀ �@U�jҴ�h������׽v��E����Of51�br	��~�l��g��/=��^3�+�N���e<�ы��˝�WCә����E;�ilD���r���l�UN���J�m�V����&�%�w7ukd�\ws.���5�[W9�&�N�*U1��%,�g/��6�����v��j�W6�EP{ ��+o��W��ޣ��T�u��W����g��͇����6�G��euka��[
�Y��&�3*{.7���#��W3��V�Q#t'ַG����I�d��(��Gt}G21��5n�Gm\�t9����A� ���e����gdMt{ݛ�gq�=��21���=�]��W��iAV+������i�^�߄��WU���?3�m�n�SU{/Q;�J�}ϱ��>�L�Ύq�����˒�
W9�qR�g�A�WN��q�d��N�O��6���fJP�mw����3��c���{F�n�Ŭw�*��^��j)�&���r��T��{]9����m(�}��>�N�󬨠�$_�N2jjݣmjꛌLd�j���mk��+�m-Յ��	xט��r��sg^j�:��-��À�5�cʜ�̿zn��	��V�n�*_$q䫰�RY�ۘVϳ:��߻8�S��ގ��5��짎F��腝�������ޘ���Fw��h�`+3
{��~4{������cj�OU�͓���*3��Ѩ�h%@�#�}�#���ΤE��_KOe�����<��W]ƴwx_i}�-���u�b*�x��i]�g�G��<�������&���w��Xw<��ov%���99���J�:�7
���D�V1[�����(�Cϵ+��:Z5%Wt��ޅ}���|��=���&�V���a,�R�{��t��㩣�(�D&�ǐ�rn��\���K'��M��[���[��+���=�z}��e��x��L��[���Zf�"K0tI�g:�8eCca��	�O�	�E7՛{0�>'���n�����w�2���d���t�I4�0�C�@-���"�9��ң.f���1�=�=衙��{���ǮFw���#��r'f;��{:w�-�ݠ�zf;\���ywy�vx>Qn���$�+Ĉ���l-�;���Fp��3q�[�j�YL�t�Uf`u������*f�.�ę3p��+�[�ɛaň�nb�>o�����><t���$CG����ܝ�*���ғ�
wc\ف;�"Ԟ}.�c��.�4�M�B_�_@�XΚ��©ߴ8�v�t�p"1�ۄ`D4Ql��32gиz���jTM�ږ���7QR|}tG�e�?YO��њ�V4Rط��+���S���7��*rQ�vcU������wt?vC�'��	������Yf��i���d*JŐE���,CwUQ�{���Q�L>�6��e{f�x��l�����(�i�;�{�b?R���3�%�(��xbWK��{}�2�7����^(�<��y'����ќ��2xs��}�t+���1���0�J0bd��E��fg��b�`��8��U��8&��yY&���R'ʺsE�伋X���޹�v�5����g�uu��v7�2�;P�Lb5�z�1�W~����G�]ЈZ_U��BnN �)��a�\)��Bk�`�H/>�80�ƞԙ�Z�����^_�
֬�p����@k+ȓ�������V�*aD�G��7���t�*3��7�a��y>��x����N���M*|!6�1�^b��%S�U׊��۶C7���;��z����7c��&�aO�j��Ԯ��]wbe+� e���c5��SE�x4��z܍��M���]�T_�:WwV�=Sd��<#�3�h�nﱫ��,�w��g,�*M����2�"}] yR̵m�R���ʒ*o2�Cn�3l0��ʿ���7��IMMQMP�������/.��H�ZKvv��vl��4����mL<ٗd���b�B�֭�����&e�X[c.c�v]�f(l�]��l�]6`�6UK�Rk�kfJ0͖�L;Bf㙉f6`�f<�t�F��v�-��ui�vܠ�Y��Sh�nf�0r�V�0�0����AfvK�K�Ў�1Y..t�ZJؙ�J�)4F�(�K\qm����k+,�J���zvH�Q�&��t���Mtۭmk��aRͿ��9�;��uo;Eڅ��V3���6-�U�gV�	i6��a�J�ja���դ��5�!F�)kT�P!� �l��-����D����'�7U _t�͓R�gIGٝ�liX��NЩ��kb�$��Ȥ��?E�5۽>a;>?%dI�4�9�eol�|�z�L����`��I��P�3*a�=��](��Jy���뒒}~[iϵ.��yV$0�=M�6������{��b7�+j�F���1|V��ޠwC|{m|�ī�{�O�M��v��7�ޒI�Z���ިe�408�o���=y���:�\���W�g��[3q�x.�r����T%w�Ub}s c�#� ����)E���z����s�Y�~������Y�[�4���,Xb?>?U?'�JO�cP�����ӻ�{��F�a�W����{g[w�7�JY�O�p-�a�Ļ���ǍEM�w�N�R�~0�X�Z�lԗEFzbr�(g_ݹ�>�U���B{�q�n�:��p�q
!8�8%4�������؂C��-���aJŔ��6Ã�
�k��P}ۀY�t��01��3�dtٜ��}9C#K3�NWj=��WT&nW�}��4E��,��fA������[yܶ����]n&�n�h�Kp�ťmrX-�
a%e.�ƚ� <I�WA��P3��+��.�[��%&[z�����=��͵�Y�l��Nr-����}^�%��FԑM������ݼ��+�e�2�;�i?��j	7�|i����[-���I8!�l��y	g+ǲvO��sgV�hC�1)�̿�Y��
���"������zs�}#w���(�V��V8���P����z}�Sʧ�����{��vť�����UF�Ê�W�������i�0�.!���*�g{�.<��I�Ȥ!kϳGv�=��=���q����O���z�{�g�>J:{���ru �:�G|�sx�N���%ˣ�{�72����+u��yx������k;�,�I!��Xl+7H0��Å�N�U*��.����,Ř��.\#�"슐�qS���NhB#6"w_
��s=b�7�U���ft��	�"�&���G���s����ŋm��O5OZ�dD��L��l�Æ
�cʾ~�6:9�(ͣ-����&?��o�б�;��w�~�r�Y�W[��F�K7�W+����E�fJ�	�f<�@��|���P'\]#��߯:QȽ:��С��E��!m�c:گ3��r�M��&�*kj7��+��r��k��8���.���K��vXQakU|�/@m�$gy_zǵ9�W������l�^�Fj-����F�q��o?i����f��ɗs�E��˻]6�Y~�֟��O�Ҙ5��B�P���l��Y
�Y�.ӱ�%�H?D���|�7�T���JS��0�ή�
pk��"޸��p�}y�f'�۷�߶c�jo٣r.˫��<Yg��=�����K�f��f�x�n�~{=j����
pY-�a4C��JuZ��U�ۮjkǪb��Ng��S-�C���by9�@��~����
!8�KXkAñJ�!&j���#M�gL�Ɩ3��[�&��VF���*��U�f�{J�lSY�b����ݼG�b�
��]�+Q&�\�6�6�t��~�eu�j�*Z��J��W8�Z��՚�l��%���j
e%���W+�)�K��ʌ��9�&����4F�R��ˑV���92��s��������y��~���q�
梑y;.�]��u�3/�7�g� �{/�@�}$(�S%�Iel(|�kS���*�@�q�m�Iߖ^پ��\.��%��[�ǰ*��	�'���o<U��˕���u&������x��?5��Grl�.�z�[�^^���~����'g��.�K��+wLe��zw��ف��%$a;�u�w�֧�W���?ZM�3|�Ak}�V̓�\I��N���Oz�I#no�g]HTwrgs�Y�;&d,=uH�Y	�P��}��������h�g<�8�1L�^7j�0L@���Z�n�n��Z�lsbKV�V���mM�]��%��ѩ��߰�	:�^5�+#����3Ӫ���e]���/vx+�2�lV=���Y�=������Ov�g�����Y<P��XT�?�2S)A���m��^��/�yB��<�ϲ�Z�:ֹ9�SB���E����7row����<�֕`d:��z�`Ȕ���k�Ӷ���8��w�)���Ы�m�mc&w"Q�|��z~�������B}�]t�rQ�GEq��w�����F�������;8z徇�Ys����߯�3]#G}�.sч�)c�����	7�H���������}~s����@��^���J����ߪ̧UU���t6[
E���!��8��7���n�s���7K���M�(]c���):;�����7S�u��Ǉwj�^I�B�N����!%S��B���N�E�d��gCY�o^@��]�}������w4Z�e�$�
����kR>T*E�=mEJ�כ���lm������!1��x�w:W����=�A�����1���]ε�Ş8nET�o@j�u�̏����<#�a������Ұ.0�ka4a�H�5�2�7B�%7B�j�S)�hp�9� �Ah[e2�e��Bch��iZ͐�/�;﯇iym��*�_��ʸJ{<�I��[p���qd�hݟt�Aݹ�)>E��6a��*�9�&eGOf�]\�]�)�.^������w�=��ǣ.�ۖ�c\!�i�OC���1Xk�.}�ɼ����5��W� 	{"F������4���c�;+��6�������b�������OJ�W��]]y,�f{7կU��6��uMU�d��K�	0�-1h�vB}�#�<b{�v�\ҁٚe��S��[S�V��rM���%�cV�꧝#"��9=-��ˌ���ʏ�Er�p�v��J�r峨��A������}}����:7~b`¸��DG=�����;�߳l�k2��p��gغ'Q��g.ۏn�^�~����U���P<Nu���g�,�v{1+�sqo��rY~DЉ�������.�'a�8����=�����;���z����#|���>̷3�������FZ��KY�[3�X2��i=Q�Fw��7>٢�T�ga�`>��s�v��}�Ǒ�t�|=�(��n�\Z���n��*����������EE��UUH�JS� UE���}G�<���R���Vw��ı� J�I�<3�o'��r\�Hy���	D!	�YT��QkL�-�-���Z���Z�T���^��	��A%� � ��(#x��� "���B
(YC\F�C��xCEU���&pqLJq���~ �"�" ��j��U�������2�F�\^{ݕS��5��a�����|��^��o�������gop���,�_K�~�_Z㤱��a��|�6�@j%�>ߗ��dn5�z�ޠ �Hp:v��<�����Cp
��@��m�� �S������]�-��.��
6腔�-��u?R9��P����
����ya�w�F��$�=�Pj�6f�%{�BC���G����;�m8�L�����Y��\�Fq(��������K�g����ߡ�޽�ǹ�E<�;�Z��Ś2#Z���m�J�;�Ƿ��*��
5x�R �F�*{��%hB�j۫��4�@3E;S�dkv<��͠)Qn���B�Ll��V���4-�Τ���� 9�X���t�1aV��ě�uk,]�L��C��1�62��y���%m|���r�3�d��A��U�@���b�	Z�o��X�,ŏ-���J�W�-֜�k��v1��e�2aҜn1���ʺ�X���P��N�ᖆ�APdQJb ��Qm`��(�@�Z*� �Q���P������h�q�q���-�S �d��A�> *�܊Q/��F{'�������S��4���0CJ�3-�����������V͏EBv�-�y0�P˟@q���+���j=e��=���#��/�nul�@w��+�ݟw?	���@A]\�H@'�������k���i�̚��;�����@Ea�PW����D�<&��RPh�Q0>Uh���x�:  +v�M�a�5�Saf8��

��F�w���>C0�3jRRQ_�,)�ے~�h�뜚Ȉd�`W�`� ~F�
�.\<�N��	�@A_��`����/�
{/��ۈ�oS��X��/���*��u);��gQ x�,W�D�;瓡Z�(+:4}���e�����%�[�+����{��.�k4�����@����Q[�XJ�A�u�.�ɉ���嬲�.��f��
ݾ���n�!�\�L����;�`j+$���p6�Sl
!mI@�b�ۤѓ�urѡ��S<� �5[uv���/��:��Sh{��#�F�K�
��CZY)P�w(�?[ꘔOI��8]?n<�!�Ӱ�1�W�W��pi�?���)����