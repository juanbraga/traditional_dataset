BZh91AY&SY~E�� I_�Px����߰����P�s�� ��-@$�&M��i���)��4ڦ�z��Ѩi�������� F�  B$E4h ��  !� hs F	�0M`�L"���G��z�����ڦ�y@  2z�skn�J��D �Dc������\V7�0ZSxO4����"k-�K6h{�s����^��6��9T�r\����N;�]˺�+vf4��y��꾓� ���D"[���T��S!EPV���b��O�,L>C��/�P�������5�j)G��J�P�I��Ah{-2��*�+��aJNs���&�����b�k]|m�~8�Ѐ��c\��2O,e���Sݞ�#�����ݖ�m��@��Ov����R-K ��{�l<'�B�> 		�� ,F,�$Ê FЁ�� BZ��c�m���$�D��]b�SX�WHy�iyj
�� [N�ⰹ���Y�!���T��t ͚rH��ʌ���5)�ٴ٦5�Ē	#���0��Ҕ��iTWl���GR���Ib�	[�!��6Yn��MZQ��� �		�&���8t�ep�S
�ZkD`A�}��=� �A ��$���+�V�G3Ye'�Ke>	2F����a�i(h�&�Ò�B���PEER��&�l�q�,�)2�كp�oK]{|]�k9����ۏy鏿S������y\P�����4ݙ`�p��//�o�&�����He�7ӳ�a��i���88��|N���k�������D =�D%�L"vbc�.Z�JU�MG��x]��|(���H䂺�ƈ,�P�w�)������=������W>�S�:>�fSu[���Y��J�� 4�cI=��dW������Q�P�0rd	��Y�B�jQ^ě��ث�-�ĐUv��=k�E��9pؘ:Ë�
18�L�z�9>|e�fz0�Q*;�i��R@rˁS��ѡy{�'m���lI
��fL6g�?�N$����,��/r���I� ?A��9�zY����h��� ����e�J�&����2Ͳ���آׄ�òc70eE�](���<&%`��Z7k;:l_��{��q�ԉ��9����P��=c�/y���0v-l�'ђR{��=}�v�+28�/ eD�ro��ki�E���a���U�^����A�<7�hM��b�H�ˋ`�#7����J�
L&�lͲ�轓��.,W�N�0۲���괢`���}�MG1�F)�Kj�ȸ�[�ҫ2�d�g땧[%œ%��M����H�
ȳR�