BZh91AY&SY5�Gv �_�Py����߰����P9� g$�ej �@!��S��@x��G��F �@z�d��J��       DM""~��4������ d @8ɓ&# &L �# C �$����&�O�i4hhh@4Ѣ��hD�%D$p'�A�1'��
�oMJ@�; 	���%�o![A���h0����ܿW�k��������;p���Ͱgkk���mE@�4)��Q�!�EK�#k8���2ܝ�+�v����ƻ��VZ��\ኔ������B�� �bpw����?�Q�	���u��V�'����`-��`�qj&y姞��JH�M˪�L̃��<��qI���ªlH��;cpb0X��ǽ���ۺ� �6��H�C�˨�d���t��۹����І�tDo:Sf���s2!oPͬ#S��f�ú"m2ĉ��ji�5H!�� К��MV� �Z�e)6Q�C�+�`Cه-�Βv}9CTӨ�dS�Z�Tπ�ᬙ�"[P�ù��Ν���Ȳ!c1ު�(-E�"nq���3�=�^�ٺcI�NEС���X�g�t���4�-,$>���j"�ʹi��h�՗�
@D2%�f�6�k&wЬkƜg�;������66�1�hA�;:�uȸ3%\�'\Zn�=�&n�;8��ᐂ?�"��f�fh
ޘ�$���:�5M]��l! O�ʷ���
O�I�of����'�]��������԰Γ��'���G��>�O+_zI!������� 4��K<�9L�̓�Aa�9��[<�#��;Je7��$@ �2����{5јͺ�Zx١l�Y7��cr�0~�7Ŏ�MLL[\29��e�����W��,�u��_>T�t|�ԝ�>��Ɂ����s$ ��6�u$\Kv��x�9��w���пp��`xyI����ث��ϳ�Ev�$XC�q�n#�˧4�� �Me�����u�;�a���m�͉��*If}%�#c�[Ȝ��N�㞨��I$f��Lyb�Y��(��5ZN#��rLBy��r�ܑ�X������&þuRF���_V��$n��R�#!��ۦ�.T`Jp��
�:аWn(��pZT�i�!P e.�k��h�c{( �����V��֍CG�Z���>\�P�1N��i�qn��YɕmH  n'.}*k`�K����9u�O�l����&�"RW�0ňs�n�q'�A�x�6?7*5�'p�u7AL�d7H��D�� ��I�����e#`Â�j&��R�s���>�F7��� D�[|_��0����*Ջ�Sn���$�����f�N^�p`:�07����rE8P�5�Gv