BZh91AY&SY��� �_�Py���������P�s���K�	T	!�M4О�5#�z���f�4��4?SI�OA0����M� �  	OQ��F�=F�h� z�=&�2i�# `F&��4� �H�4�ښ�M5=�z�(Phh�ѐ�D���P&�D�N�"��$���u��������.��C~�!A����,�t���������+2�1��J((3�sM���޽�8�*��N�-��0������R�]��%�8�U��cS�2��B�}ura��QA~Go������u�yҴ��IQ^1�i����:g��?�ͤ ��xG���A/�����s�/��۾��o�,�1�ՠ�V��h����Yc�y��w� ���*��"
���O���婄�J��#,U������,��Y2ףD>)ѐ�q���E�nJ�U�B���-�V�>�fC��b�,

)i�\�e3�ۻY��U���j���z�*f!�S������k��VdT�Cn�S̝C[�CZ];�E�<����j�(+1M�W*3�âB��ѪQ.H�X������c7Yu��$fc@�zK]B���EK�Ј,b��R����&?���!�kV�.�q��E�T���\%j���R���%:�r#%v̤A���E	5$�,5!-RI�� �AA̗�[�"]��I� ��Q���W�N�,��c{θ��#o�&��/W��qYd�ϧ�|�=�r�g��e�3��9��:�t��K��@�P >g ��
�����">�*��@�� ��+��.fZBQ�B+��-�َa:�uxs�%���&j����[��b�he�T@�9�Zy����1�n�z2&�@Ϙ��w;����Nک�6�Ϩ�ىL>�ɜ0��~w�&���!�����-�s�����6	��I3ظ�a���?ga�YK�\���^e�J��>Y��$9��L�+������x�ۚʒ&��]�(��`v��Zk.��2�q|6(��ע��� ^�4��'�BZμ�~IN|F��^v���6��<[��^�ġ�r��1A���.�l��	���%2���1Qn!')VbI�1�t��,���Y�RD3�$�*<�P�MD:������ߪ�-i u�F�e�K�EŜi.����]�5�s��ii3��ud�1cH�x�I��m4,��� u�)a2Xpf��s�`�ƬCfwfQ%)9��clp�2nݥW��L��Ӻ���P��m̬�@0/2��Ǖ&����T��N�˶l��dGV6���I`b��6��a�|
t�֘"�n=�nmu��j_�:Z]4�ү����]��BB�$k�