BZh91AY&SY��� �_�py����߰����P�p��A��	٠	"I��T�觑<D4= ��?@?I 4�  h   ��#SLA ��4d�  4d%M1 �dh��hdi�h2�$S��M!�A�0 M0�4P@3`@��@	�OrbĎ���C�q��W��H���!�B�,if�0L��sW6���X]R�3$̌2˒�QB�pQ)����-����q��J�&d�i�hfbrJ�+b�T�$�ق�SD�z����|&}̳1sg>����f������_qk�.�/"ѤP =Z�$"�/?:�D��bpa�8�v9zO�8����ֳ����R�v�ܪ~N���z:�,�g�&����L aQ�H����;.)�ǌ�	����L
�`���3N��Qr�)��a�,�rQmY
[f��l���D���q
�#B�(���D�L4�V�]@Cr��WHz��y��VY[g�hӱd���Ѣv�3�*��*�a��"X&�,����I'~�ٸ�Zƚ1�U#c!i�Ғb��#;�+p"
.p�'4rd%Dg)aS�$�G2Bź���@�+�+��Vdc��5�
�%�fHi��m��SX��a�r��RY�`�e�f�\/\�3VN�&��8�T�* 2%�xu�p����Cٙ�W6S� �1b�V2���bҞ�
6BYb�TGK[�N,]��_�Ѽt�0�r�?���Ƨ�T������s��.-�{�LA �@mɏD�-5�T�ü�M���@.��/P֚�ԣ�k�˖��2������m~��ѽ�Pd'�)]"_iA'�/E5o�Rρ���
"��dH�Xp$U^W! �l�����G0�F�'u�׏6��^��;$�mS��W%�ͩM�XE�7�D���qt����	���:�p-c�˭�j9+��:L�&z�@H�a�����}j��w�(��}+���r[:��a��0I%)H&v���B�3�e[w,�\?ui������KL��YnR[��D�Y|��W-IVjfd�aVǤ�u��! ��ڕ�� �!J��f�n����a����d��@�,T�d*I�N��BIu���W[�L2)Pȯ�bc~�iq|��2Z�B��e4w��5�}ې6�s6d�K�!p��1�\Y�a��UZzʱN*�s?��>F�����'*�j޲X'n�nxu:I']q�&YCV��G	��X�ub���J(��E�=��ƛ�Mn�- V����ٛ�C:�E2�Z)$�j/+P�6FGKN1�E�*�[�uWdHk�aZ)�$��ԋ��x�ʮ�z�j�E������e�lR��gU�0���g#�rE8P����