BZh91AY&SY��π J_�py����߰����`~}�=�J����Z
 $PS�!���zOM=I���hM P��	)��h�� �   4��d�L����L� zDJ�ɩ�OP��@ h�   �H)��H���  @hQ&��iA��ا��� h2
REE)��@$
5���0J&J"r�����L	D�DHe���"S�`��B��D!��)�
��s#����0Cm�L����M�\ѐBm4�����b�}��WI0/nYP�ט�KzWL���l����K��XL,B)�a��9�3.�Ҫh���%pg�N)�m*[��\C�5b�J�&�TxY��&�0�+⮰�gm�
Ze �eN׹5nr�2o�QE2�5�ϥUChli�����K>(���]!�qۦB��#��/A���-̉���j�`&�6 ���V�q�ʀv�Ŋ���\&BpBlji(r��	b`�+k��D�Y7L��a�SBړ�Zn�^mV��b��M�< b����;��@��9[+K�B���e,�YJ�E�� �R��"E���k|▛�N��jd$�˫��6����ү�넂�F,���U�	�T����J�o)!\׵h�`֜����{f�{V��t�z7�$��#f�6�Qw�!h�Xp�YŪDZ���-���B�B�Q���H.шf�!�e�<T��E�Qsh�f����Sv�Ţ��(�1.n����6X��Z
ϔt���m,S����T��݃iB/돨<C�l "�
���N䤁B]Y�&�IǝJ�HBs	4o`V�*��K�F"�T&CS.%�� @��8��$b`\�
1A�h�C�P�8+�(¶������Zҵ�N�����*�e�`J�2�G�v����Q ���:��?���'>	��:�Ʌ�R�B^Տ���j�����R�F-s0���Nd���C���q�$�
}�:4��?%���=�����LB�H�D��)�pAz�*.^[M��f�e3M���Jz���@X��_�1�nTۆ)2�eX��+ȴ}z�
@�R~e���ƺS�v� Ƭ誙#E�W��b�"�&@�5ü�S]I�p�aS��K`zЋH�p���^W�Ѹ"�P�d^XִFD(���˩� ���-Ǡ�<��β��p�*��,|^�q=�W���AD�N��fZ^�m�*�c7@�&�4ώ~��|7�039ls�&w��j�"7,��|�(B-3���}Z�K��w��q4�R���Hb��g%%Da���!��j��K���0,k{j%纒�R�>!�Iki��" ���5�L���[!hXe�קiD|�P��"1#�Rx�\�������,�,���0rEǤ�Q%*y�s�pV:6�nL����ÎҦ�+ƺL�և����HM�~S�h�����m�.Á0w8y)�q;�[�"$sc��`�H��q��ЉDIt�����7�ÛV���f�C����lfN�]%li`����G[�J�\��	���R�A[�M�U�5�kS��D��:GCL���Y�5�!f�5:�1���ɖQ�q,S����4��e�cM���ˏ��'s(r�9��DB�M�W�6��k���Ĵܶ^+?��H�
��� 