BZh91AY&SY�4.o _�Px���g߰����P�5� Ԃ�*	"@Ѣi�6������24z������ � 4 @   �12dф�14�&�i��&�&	��0`��$D �x�S'���yOPF��#��	 V�  H)�!	�M߼��
F�Q�|�2���ƈHW�"�^�Q��^��rr$��%�d��t2kz�KL�5�5/�BU� DK��!H�5G����T�Uj���Z��R�w����r�˨ R^bP�Ȍ�R(.nqbz�k�$ ��R$�}������@&4����� ��f�Nv<��7�r�mn�F����̦���%�,v&��؝�
�ZLR�^4F�Q��9�y�n�M�)a˞��@o!(�ޟq��T]ɣ9]{E�3�X��3���Fڏ��Zf5*j��n@4'K:���G2�IFt� ��qF�5����dv*V.6���h���˧sZaK�AF��5�N�	�d��1Ӂ�KК�<�C��B{I��V�r�dC;dx�x��;/�m��k�ռS��b4b$ѻ�-7p} .<���YH�i�.® ��j�v�&9��Ñ�<-��4w���ą+AU'(����=cL��.�J��0 � ��|��8Fy�RhQn�f_mIsP>LW]�U�B$Ɛ\�Q�ڔ�$h�0�p�shaV�M�$��bLnw����~�����-�}Jo]�?��d�4�
I �?^_;�HlFe����y�O6!�SZ�:�y5�]Lw���@.��8nVH�jy������P��Z��4�\���&D,&s1j]�X ��U��{��~߃DT������Sf����_�T [� �4)��8P���.#����bX���	ƕz�{�9<`{o�6i���@T�H�z����z�@ꔀT�uJd��g_�m]�j�c(2ny�k-&�:H��#�)�&� �,0���^7Zts��&�P$�� ��v��b�w�-k��jY���s�b�!3�:������$-��@�(+��C��PCeV�#-#,��@@�Xӿ��t�mYT�� e۠�#��ãf7�7|��'~C�M:�;OV�}7��Q	�5�vl]� ���}MV�gE�m�0�XAΜh�d��-�=}��p
�9/�U�(P�4HV�	ߔD7(h4����Ӂu���q�²�0�Ђ���?x�A���SQ4�%�K����v*k�D�2\��2��.�p�!�h\�