BZh91AY&SY�sT �_�Px����߰����P��N�b�� I2hъz&�=��Sɣ#CCA��I@ h�  �  ��H�O!2d�!�h�  �4�� �`�2��I#J6�=M� �  m#J@�c}!����b$�!>��d��DXH�H-����I#	]����:i`̏��W>��"@k�V$g�Mm����5��L��!��ԗeVWp�����l,�6SgtJ�/1r�a:�c�6\,_>���.XP�u��Y�r%���)K�T�
��6K��}���@3���Z�U�n6ѷ��܉s0����ۆ�U�Y�ZԨe��V�he[�+K'IBl�`��6� %�U:&�iҘaie����5 �FW!�$Ha4�m`.`�����!٠�b��+��%դef�k�4�KՓ�Mtj]V�T�%�S������镙&�X���3�fnX�K�x�l��w�98\!�-��A����f^���˕M]��`�=�!�9Kx�6��[�?Nە�e��ɚ�s��4�蚛4��圡A4�'OX���w�����m�I ���פ�T�95�*���vS��d�x�av�H��2� �,�f��@5�˧����9lk�@���*����{G�M-r��n�~Gpu�x���¢r٣�f<3^J$UTyw�Mi &p�:�?^��Oߛ��&8�;A�R@x�vG)V��KexU�Cb@tF�NضN'���΋%[ĥ=�������K(�X���.X�1p�z�	����7�k$���0���Z�t�K����Gj�ǃrz��7��.����A<�R�;)F�2��/� *�@�=�C��Z�+�s�J.a '�Z�����r`�W %"�)����Wj��W��4�����&u�%%�OY��4��ᨮY
�� +TM��2p�ڏ��rNj��}�)�,�r�I�|3��e�wp�a�F(�3�T:{�dA�
��d��^|�"�,�/�e'=�Mx%�8�1s��VP*��`$�r�e�؀�M�]x�Ā�%yI�~�VS�P�皐��5��z�aϜf%k$ƣY躦^�	 �a k{8�q�+CS��r�$��$塍�+F��ؠ�*P�ט�#���O���f�4����%D�hS)��"���h	�Mrk�VV��pP�DUxO9�'���e��t25=,�TT����O��UB��Tck��R@V̹�#r���Kc&KE��8��rE8P��sT