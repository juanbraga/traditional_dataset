BZh91AY&SY��U �_�py����߰����P�ѧ #	(��t	"�h M4�=M��F��@�S�$�􆆀      $D)��4�G��C�Sj ��M2dɦ�L����0Fh� 	"i5F� M�   � ��hD� �$���@��__���a#I&(�� C��HC	X����9iU�>.~��z��@�@D"��j8jk����ժ��vc6횸a�dˌ�#M9ye�攤V��tutjb<_���omM�)ip��4����;Ҩ��$HJ�ޑ	��\a��q����i$�o�=�Ֆ�)��<6�'��G#4��>j�����
YsEW2� ��'x��[3Mۈ!�	Vf��i�� L�*B �i�,ɦ�X��f�[ҖC�����8SN����hg��8g\�$4>�ͥ��=�y�� (�Ï)B#{q���]��o�c~7J� �Q$$���t �q�+[fŻ/ַ�f�� ��I"w�	2酇�`�+k%TI+��t���ij$\�����qK �̻`)�F$�K�$��Ue�n9���p���g��%�l��O٢2�����P2����2H$y[`���yxu��,:/(Ml�SfS�b&�m�.ZR>�(����wC Th�h�ic`�R�Y8u�L�Vj_-��2 -m�W+��߃M�'�4��ɑ�I�@]w:F�s��avB���VPS<�95�O�½ڿ}tUs>|��<!M3�����dw�J�����l��EsL�Y��I�Bd3$��;2~�����zM�	Nr%_���)�}t����g��N>jD���B���c����)�ŊW*I.�ܺ����hb`�� �Q���mȘ��Z�$���=SF�*�?)_��;����C������I��!R�7�k��4m7�5�	�$���*��J^�/A����|	��A'��bbmИ99IK)�"bEƝB|��'�ch�X��V��	�ߎҳ(-:�M���8��.V�Y�$�����c���[�H�I�tn2B�j�ВKsX�gF@�E
�@ZLB�����L9��	���%2����AT����ē8��n��Ҷ'Fy�I1(N�RPʆ�4 : �s��6�n��b�I�RP���X�:%�����=A��{�Y!�~��;��I�33��,i$�~� wK�Q�̷CT$��5��ظ5��Tq�:��)C���d`���Xt�4ɿ\���:
g�ؑ��/�-�@�8�e�%1yaZ��ĸ�2p��I�ԓ�AV�4ST	0���23�W"���x���#z�^���8eS2��h_j3d�d�l�Yۅ�w$S�	��uP