BZh91AY&SY��l }K߀py���������`Q  s�R��$�K>    �   ��	�$�|u�+��m輚��GmqM���S��mݝ-��첺Tu�v�k�i���4���m��N�8�CֹXVwi%EU`B��ݻ��l���[[Nv.l��q�m,� ب�sv�ˉ�$.l�]����f��A@(*�"���UF     20��j�SP24�`�#� �{&Bj��6�0���ba�eT ��12@�2 � 4JhD&Dĉ�T���C�=53��4����
H�� ��I��MP�����#S��v�s��D�E�P Q ��P
X%�����p���_�*��֯�6~��/A�M!�R*������w�;�߳��)<�� �t���	Bb�@!B� PH+BPP�JЅ(d��4IHҴ- R�B+BPJRd�(R� dR9 d�H�\�ԡ�� �҆B�@��Թ#H@�+�� R#+�.B dB��
%5.J�4!@��!@�.A���5+B� R�+�Jҹ+JҴ�J�JCHR�!�.H���)V�WR�B;z8��E���c��:S�tF[�X�ub�a�hR��&���i(��MzU�8��8��.H6"����m\����Ve7��P��1%$E�&�%�V���j1�R	J�5c��x��x��`yC.g�����(-HM⛪��Q�y��e�E
.i�2ԉ���p�8�*�˄*�KR̋X����T;�%AyG.��y5P2�`E�hP!�%���5W��62��r^I�2l:�#1%FF$KMXS1��t�:���r�骚A����q4�L�Wp�e
V(cV!Ł8b����!V<�s���W ^U|�&0�%dJ8��"I�hɨ�2J��� �n���yP-V$U���J�I�B,[#<��e
3dTKF�,�	X�Jn7
D)��},T�k �
�\�<1*����i��X+�x@������V��1B��dF�J�f�E6� �*ʀ.n��QN�*����6�������8��)���`!$ۺ�O��,�wV�\���͇U�;2O�,�x�ZqF-ҋ�vh��4Y ڪX��&rr�(.���d�\���s&n�&VX��s-HE�jnrHd
² ���yXL��������)O2혬
2Ya]P�Yx�C#����X�vY��6����wp�H.ql|)&Q�Su��(�,��)`�O��Yb�������9W�U�MY�w5P�����((,�9@���䊺�pN��tHt�I5YbhW��0"2e����d
k$WI��5�b��(��2E�&	���"`A�p���Bb s(���A�"���B�"�H�V�a�%	N�Y��nf�P����n2�B�.��U�W�����pa�b�E�ns���2�݈��7�v#$ �NN��˓',S9JD����s+�!e�0c�=$�A�!�6j��A�s
nD�@	���ܶۣk6`����u�C֏s��W˒el>�4�5��ά'�C���O"L�:s3�钅���M����a�lUWSA͕3�X��jJ��n]��gm2iz�Q6��R�dI���R�]�t�[Me�մ5�]��.�hو\M ��9���ڛMr�͎ټ�ːvq[lű�rv�:��Q�C3;]vQ�dō����B��*��ڙ;Tݕ�YXj]�ef�5s`Q�����ֶ9��-&���.+(�M����Y���t���0���L��q� E6��^���Սv�a�[�-ͭ�Q�e&4a4�Ҷn�l�Z!2Wi�V\vc.��-�Fi��T��&��(�ƚ7H�-�;(����YGaR�ׁ]�Zز�B�6&�ax���V���,�M��e�k����E����	.�!z�۫�!�[HY�KG���r�(�f���`���ftu���%�b��]�u�^ּkn��,ڒ��Cm�jku��֔6�]5͖Rۻj�[��9s�Yv���]�1%��J�7!���jnX�1.�k1�۫��SEesm� -�&������&�,�e���c,�edK���,�K]i�͊3&e�	��֤��8�K���"a	���]�� ]tm1x������k����ɉ��-�!�+ f�36��!i����L̇m�e:��/�����]5�ٶ%������v�l�ر9���Mo�Moӯި
���j��QD ���B �>H��;N���/�=a�����v�]�fVY6�d��Pb��pI��mnv�M%�̰��(��(�0�VEYaVѓj+&k1£3,�cQ�e�%�eUaDEӆV�&��(؃"*����17�k!�2s0����k5�#Y�KI�V%I�cIUK����4��a	A�d�EQR��.�c1Qj�+0�����!*�*���5'�FZ�֐�i
h�RdM	E-�CT��b�B�p��P�k1C�cD@���T�Ӵ��VRE@��
"ME��Ƞ(�HdPPj"�fE�J֤ʦZ5.����)�0���5e��6���",�Wi�6��-�(��S��c,.�0(u&IN��d�sXD��(�h6#R�d�AQ9�!�d,BU&�$(bF�ֲH���3� 2CNf�aPdьU��5�S'0�(Ժ���-e�9Z�"�!�	MR�SMo����Y@
��k=q�~�ھ��b͕�2�F�6����Bً^6�輬��������~����LR��|t�B�:�[1+\i����V3C#H�p]5�]\K������a�1vƚ0ؚ�f�(�Wk4�kjWY+Ml��bhA�����Д#@�imR�CY�e��`g\U����i�hFܦli�9LD&�lh�u��='I;��'���;R���`�ܫm���Z8�$2�m9��k\So��~��<���4%_��#���4�.�B�t�"�Ya;�fhׄ��C<�N�LFlQ��ޤ��0 AȚ @��-z�|�)�C<�!H �w"&[�%�*��=��[7g4H�~�9��U��\ϯ)Π='\2�)����t������h+ra(?kF��H�9��%f-�~�<�/G��˸d��I>����L�RѾR���J����[���"�@䝓�� xkp�5G�!vA�\LЪ ;T&�f�1��;���-t�Ȝ߽9�ލ�l由g*���~�j�zj$��&��{[=�o=Y��n�Jh;`����6�[��5)+��=�ώ{�Υ��^���H8W&��9	VX�u���}�|4�a��ۓ,�����h����vۥV�E������[z17��5~����G�j�=[��lV�a�zU`ְ�O<�9�~�c�����t���v�Ǝ��rn����h(UZW�����B�礥��@��(��*���}�Բ�U�L�,�������H��6
�q"��}�'� n5NX�,/f�*�w��Q��X��	�A��$��� �:��ث���g��T,�j���gӰ#'}�~K�I/K�ѯ6���ZR�F(3C�mv�H�z�Z�P�1�/��m��m���#Б�3gh�C���ll0��%�{X,�7i�˷]eN�������u
�s�kC6.�w��z�_���^kuFm+bט�[�7���YS5�[�7d#Ȳ�(���Op�[[H��7{]̓��~���C�?��êDҌ
r�Chm�
)J������i6(�J.��"*PɊ���$�ݽ��MKX��
\;��˸��v�� �+NfTN���'����ϖ�z9O8�q����~}�tƶ��%ǣ��
�AA5]Qv�PO�E�`�.4���ݎ��6����̃�,ɮ��+����}���k�g�g�}�왖�^����ķ��Eg���pA�Ѣ�_C�\s���]�R�_����0�ؖ�k�7��n%-��wēSU���8���Box�6��W�݁C)��p���\��5%�c��y���kv�efA<CT�(݃�ɱ�y�×�}y�,�;7���I�{�Rm%��p/�}yfLl7��BZ�V����C�M͛� �;.�_`��0�?o�G�}80�݉�Q8������4��e`"i�O;�k��"$���� �9��ޕ�5QΎ�W�����z��?w�O:�F�9��U��E���[�c��m�:��Dᎂ���<t\�1;7#!�b�����J��Rg2����S�� z��<�({���
��+ӓ�k� ��� �X-�*�z]$<�
UR<���˝�ZNQ��e�q�Ƙ�>�j/�u�bf�&�O���89�Xk���1�b(�jME$�pYF���2k���eYqU�h��E�/O��U�z}Swd!��g��Іf���W��_V9��0�ŋ������}u~�u�Q�)4ـn��j{���VZ�N�扟ؼOcah�L��@�<4
�ǣuaq��S�n�Ia��un��å&���L4���{8�j�m� ��S�t��*bw�͛����S�0
;Y{Ay��6�IG��;ޮ5h��	�1����9[C������q;�PHuu'�i��äʶ�K������M��o�B	�2�p�ȡR ��� ��S&����LV|��S�.J��.��W���Mr34N�sZZ��Y��M��ט󒻒Tc쮹�W��?>7��gTU��e���(�B�CQ*1��'�ys[���KrfəU�v�H:"��zѷ;�%���d�T��V�˼���b[��Ƃm�w:��D:��*2]P��ڸ�Vu��-SF$xK���8�V�dBg�s��3��-����320�,2:��si�Vh�k���F2�@�ۅ�W<�h��1��jŅ��@��m��ؖ��+����<�s]�h�Z��Jjhc2遹��n���,8D
<�n�p.q�ͭ��6
@�"UAl�M�ʚ�f���C�5|A5]���o���_\	��'�շ��y>б�x�t�3�妽��}��߹����8v<d��a�R/<N�|bfDvu��T���W��<��վ
����é��,��eE�1���2T]]����b�����[��l��&�����5\��Y׮��U]�Yv@U�ؚ��>��Z���e�ʱ ��Ƣ�#;�'��6�&��U?4�ǎr��o���sj�&�b����jWT%�ne:�`�:]@4�7`��a���Y���q���u��{Opj���	Ch�<m�Y����,�ET��Q۳�ٹ�ͳ���y�Wa�d��@��RAq�x����f�	ꒇ�}�HyP�/�Z�?T\
��H��� ��M��&�K�&�u�ьmmm[sD�$K<ǖOZ�&.΢�N�d��ybE�ʌY�6�3b��Q��7}�*��ʻ뙝>��Y���������`Մ!2��ߨ���u���G!����7�f�\^����W_؝M�������"�f�j��Oʅ�W�D��̠G���'y��3`L�~�^��Fw����O��7�����p�0-<����`����;x�UQ&��5�'2�	 oYNp�:�fö��%}ư�sh��r��8�7�����в_#;��+��O`9	tDК7q̓�|����CA��)�U�lO��Q���7���%t5*�`�9��/��6�Ո3�/{+��b��.����Q< b&�e���U�]-6�Ym�l��M�pj4׺�q��d��Xsnj���
�dy`��F��q��=����Op���xZ`��q28]o���_ә�u��X�f�9�Wǯ�'���1�tN+���l��C�r��މ�6�,�9��Q"���0� �_��e~�c˷<L��{{f͒�`
�!I�,>!�a(�"}���ڛ�Ҥը�st^�̹�n�	l�^�͛����15md�� N�RQwyR-��t)h6v��YDɭ٠�^��6��|y����o<f�����ӌ�hK?��_��6=��.�"Z�-��Fh��>h�,�*J�u��[�:ŧh����U�[WI|ˇga�=��My���u����T�����ט�y��)]ƍ�]i��X5[ x��^3zJ G��틛��A�m�,��Y�`龉�aۅW(� � #
	�0i���Ai��e�, �$��
-�tz�}{�P8n���:�#ºr�(�b:�eV�=~����o����豲�f�K=��L��P�Ӷ��C����z�=���r�{�ܤ�̡V�%D> ]=T&�e��]�f���{��ޡ\�m��'�メ2�e����)@��T4�m���Q���-u>B�5�w6��S�����ޭ�3 �.�Pb�`�X������g��D�d]�鬢���d����i�b)4_mY����@�Y&�
�Bd&+^����.خ�Lp�\�7� �8�*`���>SQL�7z��Xۺ�Ww��q�#���v�˧�����;Q�t�c�wS����cv={����z,��F�pE}e0��*��m�c��u�[�:��M	�\ J�FGh��76;���e��M�8Tpvf��Z�6:C�s��~eĔu�1m���C�����Ɂ��v���pf�wR��b�3T�C^��]U�gî�;Ż뎒����.���Єc����<6T����"`Y����:.�}�c��嗅G��>��IzK�jŐ�͋�ִur�~������}ڻ�=L�{�=+�=��	��6�s���]X_��r�4��x�;���>Ƣ���W>��w���+�JQx��'!�_����r+���E�D�X�d�j\���:["-�t`TTC3�-�����^d;bu1��;5�姫?���;˿����κ��a:�</�k_����T�m?B����~E�ª���l�ť5�7�ai��e�+�B(ڸVY[c1�ͨcDf+��;��+b��h�̜l�������jr
��MSYS�YG` ِ�ŷ��R���arF[e����v仮��{[3z�m�	��V���\	�H�`�������s�3Z�Z�qo�#�Mf�f".����EłZ;f,�	u�˹m*Cfk�v#B�m̓nqjQc@l������o^���fŹ�[��V��%��0�(����iAd�\gr�b?)H�L̾W#�;�e��Bˁ�՘'o�Ԑ�'�A�ǽ<q�ҩ���U�k"A1_D#j�^\u�H[H���[��y��!�xYOkگ�5�됙�
���Żښ�<�׶��B;a�G�#��nobcN�|��s,<�=ɜgex���<e6���!7�}�4bw�\V}�V"p����UU�X
3��YSts��D���g��6g;���B-)�\o�x����DǸs]`y��j<�F���s������O��^2B�!(��1�����^�����7M�'UBf�T��!�Ğ��ty4�����{s$����P�'�����6�Z��Դс��L�m���K�����RMI2�GzDF�����@�'	�x;]Xaq�7ｘr�U�Es[�BG�0��
P S��'"��R���)�s;��v�q�%��rS�5�\x8Zy[���;+[f��J����cC��ܹ���-��Q�F�� R���Ԓ�0�[kf'�>	%��٫��V3��ͦ�n�!���f���֮����J�=c�����\�E� �� �oA%�Fũ�f6�.��ٖ}>��x��[n�߶��4�\Ķ��C�CF�H�\uI��!m�[k�B�%��#0�#jЧ��N�V�&t�nr�;�E������ӹ�����v�v�
��`|�;�|z��ߟg���\�̱��m��УFd!�P�u�+�Q�_r���,I���!�k�Y�Jdw75��Țp���z*��\�K)�J˝��۫�@�`��7��Ewmj���_�Mtt]����ܶ��8mI��E�=u��s�&\��En�,���e^Ϲs_�g��y�td��Q��B�×8xmU��CsH3QqYTx�N�b�In��I�SAM&�#��3���o���~|ҙi�4����**�����?�I�k��D5R�5?&_��B�*#f�ǌ��7&��8�4]^��r��r�D�WC&*fDQ�˹���nQb�i��oU�C��\�ͦ�3C+ml��95uB`nkc&�����@���P����1��m<�~��h�o�r¡� �oX�y)�WU��Ԝ6-���tfo�h<���#0bC+&�"xD@O���nل��1��K�6�W3g�4�EK������{�4Ⱦ{��WSo&�1�#J�կe�o^�@�Fn�u{�U���2#o�[��ّ�!X���� ȅ���B0R��g!�ePM�HZd������]�3�؞ܸ��O����&d�­��-���*�W�GBf�ù�+R�O���!��{!�a$o�r*���Y=)W��掄���'}�k֬.��^��I����n���f����*�L�s�b��:�識�4�]����-��J�|�y��>WU�1�w=,w|�b6��l�G ��4��[���m�R9N�d�i�{g`�D̉�"�[�ǵ�v�z(a�4���{N��+"xڔ����q�����$�0��bR�*�ث�R"�(6_m���}�e�d=!�]г!3��v��'��r���m<��l��쳊��Ϡ���Q�ǶǛ=34-L�Q ����ղ�ZM��m5�5����t�J����eI�s����3�kC��ߵ�jz�ļ�A1|�0��U�oW�_�W����>�늢-��}�@����!\4k��]{ 9ͤT
,��k|�@�g=�0$gZ��ٻ���Z�xy���}рAp�,�����G��\������ٷ����҉�����n;�z���4`�`�#���{���V��i
&�P��e��=������mR�p��k���������C]k��v ��>�Y�B\�
}\f������|%ըc���Ä�2[(�|N�ͭ�
|:5�0��ݻ����Ñ��]lf=�g��z:�}����p	~X��?둵+��~?)9�U���f����RM�ؽ��$$sbY�����J���9V��A�&s/US�M���Z8�ޑ��:��1p�ۍF�*0�� �QH�8��0Е���wr@9'M$��{2%��J0f�f��Km���M�:��IG�e��L��ֵg3�&�7��s2)H�,�%ː���F9�ۨ��p�u�a �l���è�y�k�"���l�)��d̢�en��段�������(HMCg�?LW/z��:;i	�GV6j��ͭ2�%.B�P�m��niEu�?�.�3?��C�}.�$�
ꪮ�e�_b7ڙ�)�Y�U��?P�nLmݹS����L�K{�Ë������OZ�����B	jf<:���n���`*�=3��o��`~���C��3��J�j1�� �i�>�8��x�w����'/H�W}Wq��kJ�@��m02�骚Acg9��j#D�W6m�������@�]s��ҝmEU�_�>誉��# 7z/��5�ǷrW�ߥW��j�{˵���Z\���^�S�1�y(���'���}T �wdc�4�&��Zۇ��������|c	Y�g'�5�����,�jӖ�K�s6���'Aq���ᏐV�&��dZ�YQ�qp��y�x"�d��]��+B�w;i!�a^g�+��̿=�2W�a��t27�t*�Ѳ�E����� �a�瀻Y��O.�UU�y�65X���m�����j��F�L$_��)���WF�I�%dW{X�#�ϑI�T6��y����F��h��X7[��O��3��OH}LX��6N��f�YQ��J�SR�'4���v㞹>@Y	� ���#����spiV6��)w��56}�N몜'V������UX�l�q2���NqH���Nb�Kj`��홻
�:�s�L:;����2ar����6�~}\�12��U��z��U����	+��	U����7������cc.��t�Іe�t�\��fp<��Kq��m��L"SM(����3ע*����%ʺ �}�j]	��u�ӧ9C��d��w���Ni�n�m���{�ϗ��6����er�Lt�Mh��q'��S�����z�9��CI�Tj�~�� >�c�d�C7Q�+/�LH�^w4�PB�z�c�ewsDVI�5�Z���E��w$Ebv�!�ݸ�ؑ�9ɑs�@8s���������V�%��Sh�NZjhh�
[`�5�����ZٌU�ML8��ٙm뺻4i쳖��z�t�4�>�4�,75�s�W��V�����p�S���և���豔��-��M���BQx��96�lr��~�-]�ʑ:(O�7�t�lȗ"������:�M��##� 2�UT�ȪJ���M�ڹb{�z1��׍7XK����^�Kc��k9���C,�]G�{I>v溍��Oe���Ѥ0��(��Y3�K���s�Yf��H���ϗ�t���>o�9S�n�,��I<=Ã0�)��]*���۸��B��WM�^��U�J�B�����q��pʃVf�<W�Y�P(�gD�,�����6���P�=���</��^�3
��2��Xo<B��S�[}�J��Ѷ����{�u�Yrw���mr�P�qJz�Y��Q��퉡H�6$��o�c��H�F��n�~�0�{�(0����b����
��3�͗�{����}�Ŧ������^�#uns��Z�7�9zebPU�G�v�9A��*�`���b]x�Ǝ4sx�9��^={qI�kXVm����fm(\VԶ�CL��2�gJ�Z���`Φ�I[�3Ü�W�]��R����T�j�3�~:��wg�Y��!�|���&xT�Q������]�n�j��4҅�ށ5�}��ßM�n{�nK4�E�Þt��b����<��h5�ζ���M���O(�{���U�Fy��H��0�)Z�E���u��o6������S����MAi�X�ۡFL�. �2uN�T�]��vD�LP��� ��.��a.���ºcU�ݻ��y�a��D�)�j&���y;�:è­��ڳ�V�,;u깡ڕT�,��XN�U9���A��Ğ�N��$��4<�Z�#N0aѩ�No&��"���2�*�� A���:�m�h 4Lc�����3V�J�Iͻ!�%^=EB�(�tk>/q��7Y�@�[�j�풱B�K�c MO}KaMl����rl[�l�Z���&e�C�l0�գ.%ufKI�;�����LJ�.�fcMc-�D�uk�
��b#*��Y[��S�̱�Լ+,aqw	��c,�½�,��77�J�Mi�$��i�~��=oE�]�����Y�Q���LPj!n�n��
$f�s�?�=����}/�~/��?;�����p�~J��=�Q�v���bοUg�8ѽ=�\p�:q�p&i�ʻ�EA���e�vI�{:޹��+���C�{�$]��(�6=��)ԍ��-�軿9����޾�Umql2�P]Ō�{%�'��"�m���*-[yqnb�����-o��/=c��}]TTK������ƚV�=�YI�W2��
�y5��{'�4�og+�9�)O���DR��GWH%*��]8&�Ɂ�WCH�p�&�܊���n�o'��:���X7^���]<9�鰴܁���6e^�[ �썼��khV6X��j�����10l֖ƍ�h��v.-Mh�TC �5۽���Չz=o',5u}��g�S�be���6
��튽f��\U0�1�l�'�l3=�-lX����y��>��C�y��F�͂����Ҥ���["J���=�m�7uPt:��~�=tj|�1_�v< '	A�6{=���5�Ď�yw�ml�uM�����p�;0"��Y��[��̋/^.�&;v]ya�J�P0���e6Gi�F:��l��M��K �.���-���aj~K[�Z�7���u�\�`��/9��D�J�0��.�x�>�me>�[y���ꝼN��d��;]n�����HP�f �uᧆՋ�x���;��������ee�Z�V��t��)a���m�H� 8��[�t�R,����{m[�>�qő���F_��h׍��%�ܼ��4:.C���$福�0b�"o��<ѥr�بl��7U>�q�ϯ�[Qf�*`��	��OT;�{���\_mv�Y�^Db&�rW�ٜ�B�q�}l��u���*&>+��'�{5L��ϳu��;���e;6�)cew
�m`�7��a3
�0��=�m����"��Ȃ!�����A9�ɤ2n�F��d�F7Z�6t�tq�..L�\Κ����P�/s�ӹj.��-��6�k�u�^QlO��z��"�(	�6�]�#/ٯk�~��uw�7|�5�@k8M/[� �QG�vV)�K��u �y���]���/d*��Ѣ`T\�*^�ǌb@�����Q�q�R1'�t���:����H��q�1�0����ߧͻ�Me�U�^�ut��u[Q�.%��.�DÄn5�}||�Tۥ�c�#Xr�:�T��q�`��f��"F]���7驪��Ix��zT�l�I��┃zX�ܹ|=�N�.���.v}C=�f��k�O��R١�:�/{'��1�`�A��3�Ÿ���={��]HX�VMM8��� �l�b�i�9��s�U�/<��Xf'ӕB�l�q�}�Tpl�m���c2���1�*A9G�*��*+vh8���fq�,�>6��O�J�ke�iALB(�� ���ny+0f��;��pb�N�MQ�s^�Z��ռ)�Uac������t�~嗭:��jl0�m`;��vmuH
%�鱄V����4	5�
��@���W�x&��<;��w�r��k����dT�C��^7Z���+�蝓��+q{�q��&�8m][���t
��q�K�̨/X,�%��l8�I_��{���r߮:�1�Ҫ�E�ܞ7��n5	C8�?I3�5�1�ȍx�JmMӞ��msA�ݩ��E��]�h\T;���E�7����~��S�#�Q��q͗��*���� MT��0�Vk����Yu��3��1V\�\�v�0kJ�-��z�E�nb���"z����P��D��f����d�/��!q�J���iJ�8g�4�n�-Qt�)}nV���hX�9/Jl���p�bHH�-TRB� XG�����Y�}k�벟/Oè��χ��eߣ0���6@A�ǖi" Ny���� �:�iR�"A�R%MqֲEyyH����)�S_�ԁ�P� 2���u��TaB$N�7ҿ��)y�۶q������x~tz	 �G�uuc���?�YĶ�4w�n�(�f�v��ꊦf��]�_��7��#���g�ڦC\}��߫���+�2����h��ѣ]�tY|��6��t��/07�GO��~GX��a�U ?5�=���>���_��_���<< *+����@�2����I�{������o
>N�X�q�b�����[�H۳��"~���T ��_�?��<��#��:䇧��'*�7p��8���k�+Y��FpA�+z�u{������z������kz6�J����x�>�W���"@A�]B�J#�"�",$*��J��� �H�{!Wn;�(�n<0�ͺ�q�I�z�u7��TWrLCy0 ]O�����x����?�͜|F�����>�+��O��8}��z��W�cY����{��ÿB� nn�v��㮄���_���zr�<��n���Ī.;v�m��ܞ�(78#�YF���2{y��N�>]��EP��M2^.��w�(W�q5��׷o>}<�>���^��� ��EP����O${��`W��i0�:���0��)�=:Q^<'��Y�l�8rcP� 'y�ӣs�ߵп�� �th�q��&&z7 ���x5��4�a��s`�5�3Px�|G�� ���G������xSĊ��s�C�y�͂w�%�-Y���+�6�#w�����2��QA�|D�1=�y���%�;D������w�j�>����,EPۇev�z�K|����L�f͚���l��Dj�d>�������W[�^�Ϯ����=>r�i,�[�A�1�����l3����ਊ��p�3W����q<��A���vȱ�ӧ�/�p�X��U3r��;:� ��}~���r������|�'��y ����vL����o�o�q�����7��Ū;��{�`WW�x���ܑN$5�� 