BZh91AY&SYpE` \߀Px����߰����P>q��F9m��� �S i����4�i��ML*h� 2 5)�6PѓOS�2 2 = sbh0�2d��`�i���!�E
zԍ�(��Mf��4 h i�F���
�@%�� $�/X��"mA`���'UP!�	ȋD��}��>�Z '� J��Ph~��\yұ��0����J�`�(Q,�5i��l�!���\U]Z�B�7w4бڙ�؀��3�<�R�#X�R�c�H�o�3����w��f3�ĥ5��ٌ�ҿ-"�`q�m��4�W�M.��P��[,,$�<ϝ0[b�D���c��22� R�0��c9y*M��Ĥ��w��(W�8A�7vV�JN�j	8*�@�m�2�Ev���2
e�����3 M���YGP�5�h�᭡Ҧ�l�	à�Ż�	%�����>�Vf��^K[<�6Z˙â�����Q���e��A��Uj�Wд=P��J�GkSJZ�_�m��i �IiI ���t��߂9v	B�8��!+�B"��Hچ	#X�h2���%t"�#6� J=H�Pj�<��4��J��{Rܝ����O��o��}~uɏ�_������xyzZT@�8�j��9 ﻣ�j�Pp��=�ӏ<�?c	ҳ{�%�c4}�zηA��;Js��"]�����c�1�80J��$ɞB���}oa�z��.�����^n�hi���?ʅ0���@��nW�|D8�rU%0���j0qZ*8����~�a@�Aԁ.;�6�����D�J��� X��KaV�e�Y�o�����/��`��T�,���of��pk1�m��xYk~6�o�jI���w���\�H��$w�J�}8h�-�˳T`@%Y�0���\N���E,5\f�1�IH/G!�3J�\x�)B��`Q��p
�����Y�Q�`\<eVK���bX:e�]�����hR��-�Cjs�(,�B���sc�^��	c-�����g�II	��B!�����'�2���X�1��:/�F1�ti�D�<�x8e��ˋOFMܘbT��+D�1B%W�eC�|��Q׌��(�Ri�t��_i�C�2�u�do?\�!�i�F ��I�6�$**EL8"�$�5f(�K0����LJ�
u�2R��T�St�0f�s���J�Ȭ�yƌ���wT��`�p���3&K5���?��H�
�� 