BZh91AY&SYЧ� �߀Px����߰����P�96u��h�2tDD41&4B����y@�='��L�h1����  h   )�h���P h�@d  �0L@0	�h�h`ba"$#Sh�Sjf
mG���h4 ��h�$[�Tĉ��IX�({����E�em$p�� �����B�b
��:YFKA[W��s��qhTI�q��܎DC��*7�?-�k�׽tVW����<
�-%K���d�g �f�,�糐�]Չ����ヅ~��B��������} \;)AU��"\��CEx6�>�/�B7�y�uґ���6P����x��(���;NZ�U9IXS�=l�B���b�9�qi�hJ4,�5�{�a��V��g%��Ғm91`�VD�aMT�P�-"�5�1�Ŧ�z`�����L�u:�[7vr�gd��v���7A�+ј*��^dTz2��`�B��9F2��P$�3�Y�NF�Y"�g6��<)4:4�9��VHI�d��!'J��f,Ԙ��e`�a�V�F/��mI		.4�@�?��x	D 8�6��N�;�WuDaD#����!%6�� 50F�DJ�#���50�A���FΠ� �#,�G{�5]�'e�vL-6���_M���S�p��s�eqxy�Xb~��֮�e���[롫y����KQ���9H���_g<2�K�yHG��ck��������J�E�SCb�J�0�9�,xQRS��U〠��L�����%�gV�fH�{���˴B3{Q�7<��f����7�-�t��X:�Ŋ�g&��8*�%S�
�Xm0��,�ѐ�P�xߵ�n
�K\�@h49�
�94�-�b௪�б�"�
)�2�O����;�x+L�S��Aj�iO:�̍�U�>D�9�RUF�AÕ�B��=e]���
(
��r�iYq�*�d��g�7��=Z�JӠB3���3&����^��1����ci����0����D#��
�E�l�(�J+?s	q�E�*�i�;�N��/0B�СUٯ l*J/��8I/{��T��*0��i,�ixr����LuC�O���Lˑx�yxK�դ�h]R�d�xr�0wP��� �C;�k���f�#A��j5�s%d��C�n�-c%��𙖠���Mg���5֙CE/���:,3�0�"m�w�!�e=��ួ�d�l)��=U�$Vf%�U5�;*	��eIEE��M�E��2@"�,(W\�a~.�X�5�"B䃧9�_�j��ђ�βW+΍V��u����`�SV1�ծ,�[�a�:d�Z8`��ܑN$4)�f�