BZh91AY&SY8��= [_�Px����߰����`=�[(  qI	֐	$!��MFI��!�j26�Ѧ�H2i��� �%` ��   da�& �4d40	�10�BiMOS����@�@����& �4d40	�10�"�jzi���Q�SG� �C��PCF�D0��AQ�2B��ǝ�O�сh)� �2�yＣ��(��H ����v�5�Ҷqw]J��f4o.���p�z}�<~<���vz��s�`����d����?�˻"���K3"Pt�+��)
����T� [&��I�z�>m�P!�8q(���؜0^%���C4���<Qyg(F"���hV�d��{z֦%T���e73P6\��tE+*[��Nl�X��רφ�^P4��׺��h��x���ד�-��DG���O�xُt��.��������ʪɬ�����g�̜�o���� 8���Y��/�|}6�jٛ��7�uc���
������BƉ$��S	�>�����5��8I$���ch�L�I�q��$XWS��Q���L�9�? v�� rO9d�D�	 pa�2�����\��+(�[o�!pN�0.5�V�lu7���[��,��)뫱�]s� 6���
���F�Z��F��Ʌ:��ֳV:�;��ڢ$�mᙸ�d�̽�k���� ���tg(�A#{X�a�.�mꩉN��`j
��3S�y�̍N��Y��;�6�ka�:�[ɾ���� i$�(;	4ݹ�U95/�h�M���l�����ׁtpؓT♆��I��M����n>E��x�T^;�K�[M��T/0�c��T�����A�Z
���&�E�!�>6�4&k��31je1�|���(6K����E$�Z���ec�O�[��
�c5�CK�9����TTM̗m�t|�'�ȩ��$�5tƣ��,+sш��N����Oj�f%	%�L�4�s�M43��NF	�`�	��O%�<fc�A��k�s���N��H�	�� D%�~��2״�ٽ�lL-���0��ĵ�T1�I���VJ����Ch���U��$��R2�8���
1i"���%��${�*a����8��V�ަ0L���j7�R�n>��7u�Ͽ�����d��O��vr��|+���,D\;^��|!A����2��5���Ci��;�û��-ف���e
@:jD���:N��i�R]m�g>����[��c8/�m7�!�1��1��C2�L��$�^֭��E0N��|��a��;�R�ŋs�ey%���IƣW)�{!���	��C݄� ����+3�6��)�JM�+��0�v2p�s�"�U˱��t�Lo A4Ʊ釬���>r��0�Y��s�8?���.��!lK���ݙ8iW6\3`3$$�LL̘l1g�<���ǿ����h��ʳ[܁Bn C��<��K�����3����Z�Yw5���D�-�r�(P}?=FC�]h��
�ʊ�d�l�)���B�@hV)�`��-�GF�.�'�fF<�nQ9IË�bƇ���z'����Gষ�h.���q:������N~��q!iG��u�
 B�aX�5�ۉ�9�9\aDmd&���a:�:�V�(�@N�(�	A�MB�u1MM �BI�&���V��&0��1T�Ym�ʨǊE(dj�V��WXn/�-EG�ez0��q�0�-��j;m���q�d���z�W�]��B@���