BZh91AY&SY�٧ X_�Px����߰����`�vn� \;��$ I ����3MOP�h�4� �?@&���@ �  �   ���a2dɑ��4�# C ��D���� �    9�14L�2da0M4����$D!2�Q<�S�h&Sj<Sj��4����I F��U� ��$���@��=���Q}f�<� j||�D� H�1��;FKAf�k�3w~x��4cj!B ��8øN�gxP���^��T��ӞiK9`��s���w,Qˑa��(T#��̡�
"�	2
Jݕ����|��}ut$eL��Ǜ�~HǑ��*e5����Y��D�֙BBǷ���<	&��M'�J���^�Q	3$2ȍv1�%/SsXoA�ΒŻ������+���K,�(�h'�a��4��0\���:I�gZ0�M2C�C�$U0Q���+�"�ӕ��!�[��Ѫ%Ǚ����/.IW`�RՓ���J��Q�I��="R�Jl6W�qSkMn�lZ���!6p���i�� NN
�J�\�(3	��VY���Є�>�,��	�!믃^y��Xwy�Rbԅvt���%�o�U��2*셄�p[|3m��#
��NWM�~�8��FH�7h�H�S��7�<j���F��m᩟6e�̚�
6U�����زj���U�ē.����ds��p���!�R1���&��'�΢�T����z'&�>p�+�@�� �8>]]$�Ii0;��)���S�\�gm��ob>mY���X4(s��V�=�"̖�C�!�,��L�͕YG}"��s���{�$�b̫������F�,�]c��9� ���2�7���^,/X�Y�{>N4��~L�������V5���~��?��w�G��\�b�ӌ�s�#�! �C�N'n���+�Z��JϸYO~��J(�:������x���:K_�[v�xCx
vQ�7#�ŚcO@j�	7R�쾤PcLǿ���/�OT��
V��r�%��á��Q9����8�`�i(醈���[��H)�
���A�A�5V�$�U�iM^�Z�u m�=��ڧ��B��A��B?I��i�9�P�V��A��(T��g�ƵT�\�:�`�Z�0���05(�i*n8#Xo�BrV͛$�� ���d�d����`�!�1�Be6�7�����@��A�ԽB���r���(%>S	p�E�T'6�ƈ)ԡKؐ��|z3$��Av�N��"5Pb�U�*�)�@��(�kwń�:$	�K�R!��1*0�g1*Z�.$2%���e\2��O����6����ݴ]׈��A��s��n�+��	ۏ0@�p�s�ڹ�� �5��e�偯��R�b7����D�8���&�G���m�,9��ir��7a���ȭ8��l.Zp�U4d�j	�GD�%�����jr�eg1m3�]�EU6�HQu$B�:7�Aip�EZ�kNђ��O-�{�=����[N��2�gb�����1�� ��x�����)�(��8