BZh91AY&SY1� 3_�Px����߰����Pr�;���,�X$�	����F�h���LC���!�M2�����4CL��h%2M%?IOS�F�����@   = ���a2dɑ��4�# C �!4���G����Se=C�4=@ 4А�i���
��'�{����&,�d5�~f�?Sa�`�ѽ�h0k��8yt���։���Kg�[}exj�G[���'�z-�ID�X���$Y��.ي9���,�I$*NRGC������k���N8�Nc�R�ܘ��o��XZ�sB<`���H�;� lO&$"�k2Ს:�'2��"Q	Ԣf��g�l��z+v�!Ē^T�@����_lO��ܱr��'i�,����;���B?�f�T�j�]A̢�Vo4��+�s�PT)\jP��33ݔ{�;+�M�N��zd��[O�%���t�铰���X��^;�W��.L�w���u�<l�q���{b>�o��KA~K����}>�C��!�0���d�]oYVT@��9��8!2
�_э%�_���`ǎ�%��f#���ʂ!̨rfĹܳ@�"�P�R�&�:�f�k`U4���h(ji��P��I�A��eF��bm�������GR#�~�̬Qn�&��/�&G���}��qP�{Ӕ�թ���P�@tn���9���Ł��v	Y�4������ѦZΜg�IB�S�so���V�(��Q�Gl8�p�BZ�l�&�}A1L�+5>�M;��bL1d-�*�d�x��&{�5�P��$輂&�ɻ�9
�Ł����CW�!�2��!Y��'����C�v,%�ɕ8R��F���fdq5�,���/p�k�KR(�ba)�&���pۅt[d��0�'��QH����A$�0l�Ÿf�Xڡj=I�t�a C��r�t́�<�	P˙ЛvoB�.���PL��< o>�mSĹ�����Х0gOи�+vϨ��:���i�˦�ve�+P����A�� ��Y��H�
"X�