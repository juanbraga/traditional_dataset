BZh91AY&SYDX> �߀Px����߰����P9�d�ʩTkW@�BL��x�G��Mi��b�4i2d)4�ɀ�` LI�*d�0CL#1�M2 �A�ɓ&F�L�L$�D&��S<��z�� d0�z�!��D�D
QrDi�?W�D���a�ڢB��|m)���Eq���5 ��V��ٯG*'�"L�T>F��'�-�o0��#}nXo�;֘�v�*��L��/澗�-P��BF�s��d�4�Ww�
�5�I$M����z���<O�$Y!ɓI�y�ˊ4�7+j��T	��vW^gѥ���q � ��x3L3+"ޏAu�;�{�7�9�����T����ʒEu^^����䁔�\1�ZD�����f X�U��Z����7!�ݹ�ě���y�x4*Qôڮ��2��x�,59X��L��+���Uիk	�6"^�C���:�d�,բ�K��N,�x�pl�iQ�����H$��$@A���C���,,���"O�@�tN��#�` c�h�H$GyQ������Vx�8��sW��	��X����=Dh������������L�g׾EgmTj݆��S�G]�?�S\��]�n��N@j(q�����x)�u���h~��������a��$Q?I�9xq���^dĈ%i��U��x�~���{}b��=�����\2��N��ȇ9c��t�i=��p�e#>'���Ƨ��3���_E}�^
l"����6ρ���N�Hx���2�%g9���a<�q0�{2���zx�P.a��9�H1��ޘkzB]���Ģ������-����J㙠���ߓI[��ezɠ��i6T᪔���*�nf�&��	��*�8\/��frӀi7�H�ڢzO!�MT;�OS`�M仰�0��,�ۜ,�MF,XQ����fK�Yh�,�Y���P��Q�-r�)�a �3�Z"
K����r�����Q7�S��q9��u�W�8yq�a�$nN2q��0nW0k6���Et�ާ��	O�lu�
Q)����^UAvb����(0�hs��!�Pk�g�N�I��0(Γ$��_6π*[�
��5Lק_D�&1aB��4ҭ�j�?���:�0��bé������1K�J�"�E�=��&e�eSǳ&�N2`5W�u_�w$S�	@���