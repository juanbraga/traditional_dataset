BZh91AY&SY�Ej� �߀Py����߰����P�p:9��s����$Ry�6��F��䁞����4��#@�OU=M4i�� b i�  JhQ��P�d�i��d� @dd2d�b`ɂd ф``$ F���2��=� ��)�=hT`) �邒I�t��~$�T��2�v)�g\�����J�%0Q\X��<�g�ԃ�Y*����u��wa���B8�"�7?b���4^�i\������IhC�U�O���VT��{��1x[�� �[���?7\��d�Ɲ:�q��:�}oQ��`}<�3�$����-"C��G��y�_h��E)�b�%SÝ	�y��O�rZ"I�Ge� ,�����`�L򯆱9dh��xYfyy�={<:���			,�!8��k��	3x����8h�D.J��D\�;����h>p]&hr�&;SQ�:����E�9�"�C0���1\_�S�baDi���s��o������l�_dq�MUO�~�q�М]雓�Mx҃��9���u����OܿnJ��r	���Q^���s$�2��P̃�8�']���R{��S\2*����{��cJK�z\�݌}�ZLFfX-U�N�j�L��Pz6��-��	���{�L�M��nqd�%C��{j�a��M,S �S��.���d��e�h`��*VͰT�����!d��X�*/�Di���p�ܞR�ч6L� l&LL�Ӭl���%�4JǾ����"#�6�	"�
Z-f'Μw_N�ưB���Ly,�D���Q�*SM�|"�d���-��Y ���Vn9���򧤨L�Ȁ&L]�o�U�*D)+�e
	d��S_���PWe�ӄΘQ���emjQal2*M�4xMZ���LX¸ٷ~��șd��@�0,/2%��1wD?����f��ãX�nY�rmث&Ɠч���2��0Y��;Z��QQ�+������"�2��`޹h)1Jjn�ۨ�,��pkbl B��*"(��H^I�
DȐ��tIT��>֌!Y�H� ��d�pΌKZ̩t6,0�ۦK?š��QCPkVP�04U޷aFU��Y��:�K2�$�?\ITmaA� �kӈ��)�Z+T 