BZh91AY&SY�F� q߀Px����߰����`�5�w����š �BS
x�4���Ci6� 4ڃj4O@
Q@�    I�0h�hdb!��11	��BB&�=C!�� @�&�s F	�0M`�L$HM�z��OMI�	��b44db1@Ӫ Eؑ@	($���$�%�I�ﺦa��`H�9�͜K ���ch�2̦�f�kt���׽r���bEZSB,�Y�����Q�rd˹�ݾو됽j]b��w�n}ι,�t�*.-��y
�Z�Q/hZj����Xy^2�[��P�f�����Z����a�	y�5,0����o�@"��$$�#������R��%��9��p�P��3܏֚�@���������¸pp��p/A8e��a����	�b9�EAN�eMH��A���j�#P�Yg,=oS�$�Mn�� ]�䪉�x';G/�5��D��C̐�P��R6X5�*b�Vc�ъ��Z0�	1�F�m����j6���+C[����h��D%m6dRUmy8�D^�0L���A(�@:R��Se����0�Y�H��:HFjI0Q��É)���b��RY������+ͫa�����CmL�!�M]#wQ6���C1lL� �g�@�C��816�m=*Rr�������dDAX�a� Sf�*�*�]�!�I��m�hH\��b�����][+��&L�wd�c	dP��F�S��iY �.˰(?�(�3�]ݷڒ�!4̢�g�fU��S��� I�fg�P|=��$Bi,��$�@$g|����|�) 8���n�1%I�V�?z#`	N��'y.Ɏm]�$���)q���g3��C������p/V�N3��3Ē䊅���҅��9��⹴�iK�s�8 .�п%���� �q؏���:�,d�K�I�O^����a1׹�{�V�
-[�K2�Of��u� ���/k�B ����
v#D������з�,���RD���a ��q�2�%�:
�2�@ݗ��Ydg�ġ��I
�M�^H���?.t���$$���2K%
w����sƄE�?5���$�:/�P\g��I!�S�z�?2�l��Y�@��m1��y��'���J}�&n:,j��� H{� ���i�b�W��L3&I8�%�,��V��4A�N�fĄPo�����(�t����'�Qp]��Y9u�L�
�Ǒ�a"���g�0���R�sA�H^^%R�ᴡ�)'����J^T��:�x��X�6�OO(�U{ Ąt�G��_60HV��2N�v�.�� �*EOл,�����]�J�j�}1)DJa7���2��:ڶEU�&����'��`�o����C6w0H.i!;�N�eh�����L��WL���b٠>�i 	��H�]���
���=�%������܍c�0��<�:�Y��)�u� �i�ߣ���[�.�p�!���