BZh91AY&SYMLO� �_�px����߰����P�8� pΪ"�Wl	$&�'���&��b=M��M hO@&����F�     $$$
yC!�2@   dhs F	�0M`�L"RhA4d�Bf����4��OQQ ���R�@h � B����{�]}v�A�w
��{����!��BD�
�"G��8=X� �0.����#?G�a���n<�	�ʆq�p���ΪU�;Z�e��!R6�-#�2tʗ?����2n�X��8��D5�{��� Ԭ�U�v�i��w:���Ldc&͛M�;��i!�nV�'b�]����c��#L6������eE��v��� �*h�R��C�| �`-:lw6ئĐ22���(�p)�2��H�Z.��B<!֓AV$h��)Z`��
�2��%U��*�9p�5n��V�����J��g[�%�C Ud!�TL#a�e��H�!���D@�
Z��PD]Z+ܲ�2_&�퉄��9���$�AjU,��"Q��-�&�f�0��F�gv˖Xڐ"+B �v�LĩNīl�$E��<��Xz
����M�������I�����U�B��,`�zߖ�2ϋ
�FM+L��m�FBs�(k�ц�2d	&�f�;��]��ukވlZ�q��9z��jx�u�7J�A���:���tv|��+>�S��x�D]S��:�X��N�ۇ� 54������3��x�\ w@|�h���:��Yg0V��U�)'.�qL�6�u��O�=U��w����O�U�d�[�#f�� �p���)G4WN����`'�C$�c�J[���Tyr4�@���U؃��3Hʴk��<��,Ɯf#`�O�
�aw�Ҭ'9O"�!��)��^]�˘�-u�J�^ �spm��P�U��h�����	m������Lw=I��[��./���Pōzp��F�h�x��FVfL5��t5���#����V8,6=�6Ip<f��A�\xyB���BZPs5k�*���X��8"��d	d�|�)8��.���r�)2��V%5�x��IQ*�/F�5��qWx�.��(А��&臇B�@�YS�U�/���+ ca��ηY*��8E�ad���4;A���-�Q8��4l���U���I
�(4�^���u�N�����H�d����7��Ѩ�|e��g�-2L��b��{���%Up����2"�P��(���8���Z�fU��0��ՂSf[˕�fٺf�@̙��e�#�.�p� ����