BZh91AY&SYF �� �߀Px����߰����Pp�QDی���%�$�4hM2b�G��4i�Ѧ���a4�	�H�H� mCM   %=D��@Sh��  M ���a2dɑ��4�# C �!ҧ�G���#ڞ�yM �Q�zOS"���"� ���� (Y�w�����e<@X�yA�p@�A��r%�������_f���El�R
��2I3+&یħ�d�7W��'��i'���[��KXj�L	0��X,����L�_�б��7�6(M�ޔg���9(�[t.[q���S�F�T��e��&��u����}�� D,0i]�wNx��ķ���e;ҁ&��S�λ7q��]�mY�Sb��h$���Ʌ�JZZ�%RF�{і&�KF�q@RRX����MHb�ZM$kbuL]��q��4W����Uʕ����f2�h�w�̨�b*����;�q`��`oW.Φ@<����g1t��%�)��V*�29��$���My�4հcM[�Uh����Y���ʊI$�G0X�[�r���Q+�p�L)7��-kc\��ᩝ�^�B�w�^�D)jl��uY7U�':0P�#7�b)���p�����H��UT�D��h���#���0�c�UǏV)gu�L�!L����l�!f�B���(��0�!� ������u�U2D�0R7�@���4���/��(����A�6W��5�wX�2ѽ��<y}!&~��o�^=��I��<�#Mu8��8��?�Ё �8�yϽ���Nq�&@�Դ0��`�3oŃ�z�D��� ��H�����|S�{ӹ.���������*���#�C����t�I�}�.��=��=b�1k'N/ARz�YJza=ƌ�N͍c��`')����[�(�I^�į�{�r�T����5�R8���"��L�5X�z/��Y�&Z&Gi����L�@���\71�d���P� ��j�WDjbP�yNI�p�Gs�]�Ƀ�r���Ex��Rrρ�$#Ղ������~Bq��NZh�]���S�Vȫ�=��h*KXfL5�g��l�s�ϔ%�c��7ڑ| /����u'T9���u᱅As��#�Z�+}Q*�д8-P�ri�gA`;L-둱R������CE�a�V���
dա�f�A��I h��l�Cpf�� ��d�sj�@�j�E<R���9�ȗv:��@���m9���ڮd�G3���胪�� ��O*=�-)9����t���b�]�I����w�n]͙��(F�	��y,�F�݁��O�T�&�x:X�D�AGX�Y6���d��� "XP�*���j�R�ҍ��5���ٳ9:8lo�p0PY6� �*��b՝c%�a��D�T����M79o��dm/P������#1����2rr��ܑN$�=o�