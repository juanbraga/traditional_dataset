BZh91AY&SYD�� _�Py����߰����`|���1�X�2BIL�&)���#DɁ��	���S� ��x��     OMDz���@ �@  BDSF���z�24@�dɦ�L����0Fh� 	�6��z0��4ޔh�4i�=E$���Av$R��b�����'e��e��H�H�è����I��1�x2l�ASV5�����87�$4��G�6n��Ҍ�H�r��mL֢�BX��M$�*8 �BA�EA�ל˻YD���P���bQ/ˈ| �c!ˋ��oZ�Ǔ�u�Hc���2늰�� 3���\��I c1�B�8Y��|l�i 6�3�r��J�?K˳i,q��gCSo�Q>��ʃ�-���щ4ҳD0V��i�Q����9W�� �("h�ʝ	�D(��@�XjaZ4�I��Ă1ʻD��Vs�K uل�͏,�Z1�AL><���%U� �V�V^K^��=�;r��f�C`��i�\�d4��jȧp�{*�YBf�)EɵgmM�$*jF�������UfEN$���\����4��DFT����!g, ��h62�#G+2���˓��Β&�ۉ�Q�X�dN\��@zb4�.���km�%Y�rf���c(��û�dQ?�y����p�rH$|���������+|�&&��ulo\�2��%�-b��24h1��}F,��mT����� l��E1.�]e�v���^��X�9_8Ѐ���5#O��_�����˘5j�7�.�����y2L�n���JM��J��3��I�%ElK��^GjF�o�Tb@j	��.��?A�Zh7��T���B�<+��y%ތB���J.�ae7���,ڈ�U�JXf�at������i%ս���s�xIUW�T�ܮx��r�� i��?C8��6Z���I�M�S@���N~6���Sb	���S�Z43��]s	�2!�`�p����9 �H���4�>��D�'JY"��?�@�r;K�ɜEII9^��hMXz�μPY�k�e���g&T/����wB>PS��M�(o$��
V#}^�ȳgHcQ9����)�=|����kd"e1:�Ϛ�U���| �Rca�0�f�'��qO鬉xʪ�ّ��X�<� �v.�h�b������ard�Q�%��:�h�OKlcDA$�L��	���OoV�@pJ�mRp�wA��B�.�����X)L�x�F@D\Z�n��6&�b�;���㨡�
q�r�MA���8{�5����W�D=��d6�[A��q;�%\�� {.ޅ�d�#��l\P8HT객g��Y�=��K�)^V���ٷ�&�0�����tK
m,j����UfTE�b�t�T�O���P����@�L�e�lz�00E�@O4
�wO�W]EL�VdBr6"�=�1{���X}FJ��Ʀ���d�r�,��Z���d�m������MZ���`����"�(H"r�d 