BZh91AY&SY��� ?_�Px����߰����   P]�1�;����IL�&��b�Si=O4&�SMD��S�S�m1 ф h" �z��6�~�MF��@  �2d�L&F@��M#4i��OD��=OD���yC�z@���CM���D� Q� x(��s���KJ����k����X�m.悬�m6��7ElC���\�XX�M#����8���$na
J�����X���Q��(eN�J_�dBT�˒A�6�P�v�f��]�6�o^��شڪ~��<�y].g�߂8sv	�kQh_^b�@�J50�<�[L�ʃ��Ѩ.��ONS�6�(]^s[llm�[m�NN�<��J\<�,T�;Rl�>[)����^iA�lg�H=U%eY��Nv�Y���5c"����;�c�4{I,�Y*޴D��:��?m��>]��'+�4�ͧ�)+O�/��P0�;�9�2��Œ�h��_ K wN��6���0�QJ�c��!{���f8p�<%7�)X�2�T�@H����J�2�.��t���&f^-�c�eV�!Tըz�$�SF�BC�+;�7���
��"�=N���=l�<F��	ʅ6��!�l.�Tk2�	h�i��_�*Sa�*ex��X���K�W6%;�g�A]�z�L���HkN���j����r��a�6a��ǄbU�FQ�패D|%���
�H�l}U2�\L�Z��i�Bs4�sgXn-5�B��\Fi�����xh9��P�iS�%=��T�A(_���\�)Y"N=p�T�{7-)�Et�n"C�!uvl���a+�ԛ
R���"���Lq^�8R�q�m�0iT�8%��a�d�%�19\j(���_y,f���$�Q��J��J�s2�	���y���㙃ˀ�D�a��HƎ�X���ʦ9=U.�I�z���'=�4��>@�6�JzBC�	N��@`[�Yn$��U9���יִ�l1(��SC �ɐ[7�	�����"�(H��Ӏ