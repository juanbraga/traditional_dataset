BZh91AY&SYh/d ��߀py���g߰����`��|�7
T�	aj� UY�        �����     
@@�(F���#U��-tJ�M����um��K6��n��Ƹ��.b��w.\M[dѦ��P  � n�l�� P�Cd�J�J�&������EM 0& C���Z��4��L�1dH*���D�� "� �F���  �����,�� S��(JH�dPP0�*�4)
  �@
c ���Ŧ�U*� bi@ A� �w����"
� %J�4�@Fhѓ�F"����*�h F� �h�L�1�2`� 4a��T�*J4�2i�  &�`�$4 jj~�A��!�F�j0�&�R����4h�   4�cŷd�bE2Δ���Ҹ�" ��{�TZ�UM@���� DAZ	���HA�4�DD$���H�����j��?��$ؒx�X�l��wg�L��Uv� R! XBH�� ���@X� @�� , ,$�P"�"�E $�,	 �BE��E$�d $�E��$�)T�) R@��H �@�Ed,��uw��L
5��	S�nz�;�DD' ;_�)_�@��d\�_Ji�����N�CIv���b�-Nev�
5�h�+E��ɛ4ѷ�+�ǯ^Eh=?��1�n��>j�/��V^ܡ+�n�2����h��]ۦ��!e0�!!r��O.%��n�HٻY -J���6��m5Y:�m�1S̏*G�k4��aZ�!��-	X�SL�,.n������P�[e�`�.�4���n�}�e}4�u/%31-E7n!�}��SEMxE�&��H�qS0qd��A�$�˲u�k̒�� b7������NJۖɂaR&P��;R�ɺ��v�tҭ��HL�Dj�,kɘ�.Z�ޚ�X@6�m��QӶ��+�Gd��d��$-����WL?͗0˵�&�t�"�z)n�⥩�&�&��)=�SmPE������K�k74c2�Z�C/-�.�I^�w�T�x����k�bPVq��4X��蘥MYˈ�q�6�c�GQ� ��ت�1��ˈn	��X�yni6f�[.�~�n9�j��k,圸b�@x�,D̶�L E
�2e�&��%p,�E7�x���Ҽ?���t޳�o�=��2,0�I<a�<`Quh��uh(������"�m�V*���X���b�,W{��Xc�_9ۇV�+R��.���ƭ�mQv� !���R���i�p��[��JD��ni�G%k�u�̽,����%]�l���/
�L3u� � �OJ�FTKM*ɇZ�!�6[�T���w��R��R�l��יe	�a�y�D�0��42]�?T�.' [��B ��pT�W�N<C'w��-����2
!쉨%9��)QP���ˤ�Ȥ�MÕbhŶQb�+K�z6ݸNy32.� ��np8 Rq���99�+b��u0޸&Q8\`V�Q4]�.)����,S��Q���1�ՙp�$L��{��C��o�����I�+��Z˂h,��7�PfCqPm�֓R�2��z4[��fV�OSo&�-he��E�vwx��4&��d�m2�r�w�:�\I���dt�j٣��b�V��)
P;�M�۩a�m��ws^�	�mI[ڽ��G5˫�<����̚%C�'Y<佷Y�rȈ���d�T����e h]F�����櫧�Xt���S��H��&E� �d�NW���
0)&�ݒ� Bպ���[e�k��h��(�q0��)T��圁�%�/"��/v�<�]V�ii+�À���`JF[k$�f�1cDd�.�ʪ\4����e�0T*PT���f��Sa�!�P�2��Cf�M�u۽��b���v�L�Z9ZX� (�5I����]f�չ� �!bò�S/RvB۫eVfɈ��a97��A%h[6<x�h��CA�e���6��`9D�ܦ/?j��j��BSĕ���6+n�ɚmB�*w������=�T��sMA�U��oj�+�k����#0���Df;$�"Q�Ю�8(H���.,���H��Z��k)��ZE���ۢ�f%c&I �i�KHL��U�;�e´klQ{��v�`��W+fB�wf��6��	[&�����F���6�V^�2��f�p\,�BCp�@Ƙ��؋'�,:o������Y�������|���1;�N�?g��,B���5�~K��A���?l�y��^���iR��Һض� ��m6�rl�$�udm�"�[{a3P2C���1h̚��J�e���X�X����z��Y����\hh^#���{cM�R;�Zk����ZJ��a�[3f/9tt	��Ëm�q��5���d�c��c�����T������[iJX�D5.�iM�f��^�([�kH�퍵Bf.m���]�J���j�kn[Y�ؚ.���u�]U��k�v����%���КVl�-6�7ɋ������>Y�\S�VgJ�#��� ��e�l��F� e*=yj3]vn����:1�I�v�������+�3�vn5������#�,54�Ҕ�;^�pܦ5mԸ�v���k2�����@�h]�u��T��)��iX��`���5�E���EF���&���\�!-*�kAqУ�i�S]�\S;dʚ6۴ݙR�l[�q�)]ԋ܋f!g8�]���hD�Kl�2���VZI�CBe�4CM�5���˯[�����k�ZVc˵����ۈʦZ��2��ז���5&%vu��밵����][+�6ڌ�Yf�*�`�n�������\��]Z^�\�]��k,�r� ���I��#6�.�ceH�,�Z`��e�n�u&�g+V�v�4Wkk����.6W3,%�a��%���m�g��x���F\�&��il��7q�\��K�7Z�&Z��l�k��:Va�E��T��i�al�4vBc$W��d���;��ckn��	a��<�L@
m��I��.-��j��*@Z[`�׉J��a׋mn����&��!SM�;gR+un-��R[i���Y��f�i��u�d�&�WX���@%���9����#��am����ƛh�*@]k�ֲ�c"�UkEU�^ڽ`���g�#�/6ٶ<TsGfih�z����[�GA�:;b�aV\�!e�-M�7�.f���sV�˦!)��v�m��[k���1��2�2�sv���mbMͥ�%���K sKp�7[fD�*�u��,bbm�l1���b�5�CSA*��/k���z�l޼��r�K��i��cgL�-�ٵ�ֺ���Ĺp�
Z��B�5+Eрkq�k��4"#tuάv�P��7_%�VU��m��W�l��ٚ7Қ0mtԷ0Y��"�W��W0�{J�5������*KM��m�5��h�QY6ֵ�k��f�1t��tN��mm�b��B��#K5f�4�91t���ZB�-�:��~.i��� $����4N�y�۱A�,,9��D�ϗ��DT�G�|�$��� ����`H� ~�'Cl��@+!�I2O�I6�<H,4���HT�=B�=N$Y4�<C�$6�bH,�	4����'^><Lea<�2&��,�_}�m�6ì�3��(q�C7E1�z���9�0�oF_mU-3�U�UX�	�3 �A�ó��VK�%jܺ�`�5�N�%��q�3 ����\�O۵�{,ͤ����Ztn��wֺU�����jqJ��X"S�u,P	��:0|.���������S"CD5��e��fّj�x�c��ɶ��շ�j�K2E݇LeԆ�m�p+�A�*4�Ju�m�:��{�#[c2��^f��%�Y���d3�5|����Υ�g�����D�  ��xo�~�#Nkx���v�ە �s��sf������Jz�蚙��J�J�ٰ5��U��K��\�8��EX�M�hY�7Q%ՆZ$;��2%ˬ��*K��%hi��j���K����&�Q�;�q����`�(i��^�4����õ����"huvvV�6\[y��B��M�f5�X��K�<��n�D9��#�\]X��f٣p��\��qζ����^���F�Z�۫�Ն�u����3v���i���2в�n\�D�T�9���s(��`�8�ƣ5�ڐ���N�;�N�Ԇi�R���{jV̛lm��(�Q�#�E��(�RZgI��6\;mr��^� �a���0m<�zN��@�E�(BE�����%`
���F�`@yܒHghC=̪����z�
����h��X�#"�TX1AQDQTUAX��V(�&���5J��(*���1�U����E���* �"�<�5��h�T��*�1��]Z��Q��0QA�������1EDF	+
����o�8��DP`�X��*��EݱEPT��X�X��EEDV)���Y�X�#��EAVDEDX���7j*�_l�}J#8�������DE^P���U�-¦YQ�b��V=j�*�Q���/2�������5TV1#DV,�A���aE�R�:!]�U��E��1��"*#��;jLlb+��*XS����YYPO�"���B���4AT�H���#�Ԭ�b���H�ը�`�kv�/8,EU��U*���SM�(�(�"(���X��X�UE�Z�U�U��iオ"���7j,EEV(���s�s�h� ��7,�V,���M}绦�Q���C�[j���S�UU�U�(�~��v͢*1F"�*��ȣ���b��DX������	�[�c#�� qv{<�=+CaB�hZ�g�o��n���;f"(�핊yeT�W�QA����t�Z?s��1U�m��]}r+���w�� �%H��EQ2�ݓ^��uv`UTc��U�O
�ٺ��۬��[y8�`�u��H�YLeA;����/�U�J��,X��%����"oۆSYV%J/;�iN��Wu����QG�\j�*(��b�ڲ`��*�<��x�E|��y���>����X���+��R�y][���痻Ѓ����ֵ�=�`���c�(���T]��Q���er�0QM}��t�������o4'�A8�� ̣��k﹯��q�Q�L�)3��SԠ�ZϚ�Կ� p}���O���ޑŖ8Aj��;_-��q
��E,�w7n&e療�y�=M�w�貨ʆ��R����vN(1�)�nE�}��{�QYR�u�=���Q�p��+AE�PG>l1��ዉ��'|�>4l��xʒ��@!�@:���z���|�}?/��\�뻻�7�|+w�y>F33�<���"��Q\O~;χg\�N�j�����W�D{|pY�S7s��M��ˉY�9�b���[�uz�^�*�Ki���۱X�^wG�f�4�h�����1-,�kZSm�+Z�M۷L�/2�,���g��|�![kJ6�S[r��{ IN�0~�"����Y��Qg]��®s�o���v�ƈ��5���yl^���{X��D��
���ёM�|��J�5fXQe-Ք�.&�}O����m�rэ{�Xӗ;�֑X(_p����e]�V���iU��s�[M=��c�����Ǧ�0� q^��Ec�#> �¢�N��^ק<u��/�}|�s_b"�R�����|��y"�-���"�w���~2�{Otw�S=�9�	��_�-���>�\��
��X�tj��eb�=I���#��Z���F��������aآ�w��>�������kS�Z/��T��y��~����Ě�����TX�� �Z���
�3����sY8^�1a�5��/O�"�(r����>���W� �
j�k㎙Ԙ��K���ƜE�c�1���̱ CT�����-��uN�b�2��b`�1�<�߽��Y�MH]�}E���c
��$a0J��n\�\\f`��
D����]HXiZXK
8�*�T��ٖ�Kobiui�m!�q+W&����%n��$�ىpM���$yB��b ~�Nn��h���%� �R?{;-�D�Dq�̡8�!���\Ӏ ab�-d*o<<k�J�2�f�q+�^q���0� I�p�u]�.1��,��R��c����T8�.��x�I6_~�1 H�?b��C����E}�(�>��O;���~|��!��F�����uX����[W��ړL��k��('�D�����MN��&��Nڐ�05�̓9c��$�q�~U���4�C��4��8�/,
�lY ��_�W���o�r��F�!��M���EDX�& ���ɣV�La�S��0F)n$#�~A��rz��uI}ho�2�hi�N��So;_=�lE8�}�4�NU � ��Ғ":�5�R8$��a�gB�^��7ix��1�Jq�1�������|�A .ܹKj�J���#V Tiz��i�}�X6���"r�1�(�(�NП����,(�
�_)�D(ȹ�Փ��昙���n	ٖLY�>��aٲ�����Fe/��D�pa��#a������8DnM�
��"<X>�eĳ����}�c���Yf5�z`�L��
 �e��q�6�6& ��9QZ\?�������_GvʹH�& ����7&$[?DX�`��x��Ɯ�e��X�"(X4G롌X��`47MXb{]4}B2\�
�0��M��	pH4�11��q�k��b��DT��=t�~U
|MAk%���(��F�P!Wږ��!��,��L$�)8�R�z��1j�P$'�\�,ӡ�ƫ���f҅�!��)�qn�'Y����pD�!�� 6�C@�g�'�����ҏ�<~��9K���g��g����U���]��j.��c���D��8h�L	:�H�/�3s�~"-5�����%�Z�G�9>�J��P�k,X*�i��e�{$�GZ�ٶ�lĺ�)��JK��ib�=��M��U-��X皎.��r���ߛ�cm��:S���I�10���[Fz�G[Gv�vH҇�o�:��Y����rrLU�A]?�����"_<��Qk�>`�1��ff����k�	n�a�(��x0�G�1�\�#K��-��@ٓB4U��Do�v����J-�-�0 "�˃0��b�A�׆I�X��0ά����c�l����J���J�Q��4�>�* ���A�`
�j�X��&c#L���q��
8P�*�dl����	�5´V�J4�h�j��K�BWc�D�M��u\�]��j%�\�9 ����ȇ���%��i��7� RH�O��,oݢm�c�ZX�8�7�[o�h5Z��$a��͘�� E���,+kd�qtG�~��ܮ��E�Z{�B�q�d]�(M�oRK��se:<�ޗ�5ϻ+U�q#�Jbt��bT���Ҷw���t��d ��4w]�
��$����k�΅g<
�֕���Dҍ��q����6�O�M�P�*r���t�&s��G\���lT6�c#J�6)�6�����y��;�~���$��:Q�վ�~PҰ��P�h P2}[zs  z�n2�����r��.ceN2���rF7k��� 8�hה��	&��#����x{^QD��1b&��J{���O���,	�q�����l���F�������<  8��I'&m���B!��R@m� L��`Ǐ_33�F�#�MyӋ�������Қ����P�ֈ�s2���Dy4=�"����6>�@��Se�ڏ��j��ǂ�y��_��e�t�f=���wUY��l�8��D{Uk]R���[���ė�(ӗ�$G�����T��T;蟇�"LM� x��n�� �&�̈+�י���}k��ꧩ��C]�b��O?>C����#}X�#�F�꯹����*N
~�N�D��,��� �����0B�9G/Fyyo��(�������3���(~;t=j� @�>�F��B� ������Z*g_�>v�����埛7��F��<I�(��3�� 0��eNBW
�d@�L�s&�vX�2�P"@�����8|� 		���?a+ �ٙ�5D.~~R���ϙ�z�8���7�f(,�&�� ��1g7�Z�|yh��˲��yr���f��w��h����,5!���.�Ƭtŉ��f���kKBZ���6��f�S9�,�Ѷ�niv]]qk��.W{��B5�N�EE��H�x@��D��s�x���l�EUm5�7�6O�J��)���[Jb�~�@6�Ŋ G��v7OW�t<�1�����=f�]K�}���@�|b�|~�1<��!�]�3 I?M������ȑ�H��L��E�&X�@;&�Q�� D`�_�ܘ���ŉ6E(�8A$�+��#	�L��"l0�  /������Ҩ�b���Ã�:RkJ����'�7I|�,Gğ�\w���TD��
s��^��gA�Y^����O�)�/����PҫP�}j�Tn��T�ʋ�w�u���++x��\2���M����LW��u�^?�wK�$�;�L
0[�8�=�"D1�{�3v��-'�]:��~\�q��ݤ�����m߶w��[���O���	[~�=��y�� o"[mָZ�޽�>���?l��M���)���/h�|,D\�{���?a�sZ��/z�pf�J���4kt;�;8�:XlG�n��#|X�1� F��-u� �w��X)U�E6�Ӯ�����!��B� ���΅�!�ʹ��=LmTMj���v�n��o�Wv���9�;�k���4��^*�2�w��;E�O�ʣ0  jO�z�~~|��>��Բ��#B�L�}χ��?,� T��O=y����W���UQ��.��y|~޲�{�<k�b�s0տ�\��j&���|f�_��5/.���~y���f����e�W�K=kz˦�[;BVφ���sds��Jj"0�v۰h�b  0�|A!+��1~�.�������p)�5�,
�jZ������ww�y�����U#�9��{j�|��|�����頍H*��^�hۢ
��R�s��U�{��Y�~~n�f$��֚	a&,Ͽ;������N8b�`{n�" i1�0��l۱*c���4��}���9�y�<��ÿ�l>��u+s3��}���׶���P�^HG����A��}!-�/��|�-54Ǯ�qP��	V�Q�7�$�/�RQr�����ե���ׯ୚�k>��� �@T���2�0H$$]��E+	y,�2R�UƂ]��2f�Z٥�{Vk�m�%<�}G����Z��eٕ�r�W�u�R�͈���!� 򊇬���X��[��~�P���"����S�~8Q"���ſ�:��[���Q�"d�>1Vb�Ӭ�?B��UytI�RR룝W�Pq������৾����U`�V��]���?-k2>,ңy��d�L���4�E�(�Kϱ��=N�`����r�,#�H��)PU����DK�ts�v�;r�D�f��!�-��%KQCEH��M�*�q,���Ɠ̦mC��B���f��<�n,��DM�g������ٙL*?�al�c�p�T]�t>"(��6�����"�f��Tj Vvo��HEL_�1�K��(�EA&9à��e`8��P2} �i�*�p��A>��r��Ho � K�b�8�L���M��N�d�yn((<�c�fX�-k����'��g��᝹ΎQ|f��dEp�3�P�O���������g�g�b���{�hƈ�v�ه�:"c�娌�`mi��g���2�.*�ڷsdAu�w׸�<u�Y2.�½M��s�ʠ7A_;��*l�+���<��t4�1�p���
ge9�����p�,���^{+lˏ5��(��`KR"����Nf�&Х��LS3!q�"&��XS�ԕ�kK�@0�ɖ��O��F�<E!���3|�I�:�I2��T�+�;��y��X3�т�o$v��:EcU��*���0v˂裂����Ewot��vv<�{�$���ĭ���շ��p�-��ڐ���g5�C�d�ɳm�R�a:V�)gQ��nޭ#��;j��޻T���������v�[X3��m�r\���fum:gU�q7�Vk�e�5�F��zG�1�:�=�P��2���O#��#��:&�3�P�2�D.Mm��v�u�Jh��&��L2�{@�ĺ[t	��V�������@-��i��ɶ�-X�a��A�cZ8����W��u;-�]4��E��f�Yq�]���6��(K���vqH�jW8oP.1fճaUS�l�]����g��v��Վ�U�ɻ&Еe�˩�g�`l���V�W�J�S���v08�\�/b�Ŏ�i�F��ˀj��s�ˍmٺ7tjW%
TE�l�!dd��We�����wM����ݼi��
��fۚM��n2p�&�p�
D�4��YI�t#I�:j�i�fuQW�>%�F����M�*3��:��֯�%֝��w��u���Vw܏ik���?eȝ}3�7��s�ǳ
�Fwg	1]��U��_u�4q_���̀,Z����9�� r�ഭe�:�V�D��
��Gtp���H��8H8(�i���F����;;�Sc�2\&Lt�(��e-ˍ5����Q]�����g���(�Q>�zˡ<!��$�Li�e1���JU&~P����s�e�9-p�+]�k�>B�G
V�ָB=`���/{O]��O���붯��}����1Ee�__����။�V��4g�n��Bn���!i��ی�ߣ���v��ּ+�f����TFO��Mߛ�9��Z�x��e���i)[���*	��%3��#d�W������\��Auk�D�o�����c�<ceU�TZ�j�ϸN*��s}��Cu��ҳ���K�#���SQ�1BA��xl}}y?L3����zg۱�ڎ!処>���v�eA�[����t����{�Gм�����?wW�Ԥ4�$��
>a'�_m��~[Qr)�R[��^ߺ!̹3iC`"���r�5�6���@�XP7.��_W��v�jUg�0G��j�7х]���Mw�b�������J`��k�1�^��^�`�yQ���HDߺ�1��"Ϭ"��|}�O�x��"owjm3j�	pԃ�v�ɣ���ĹKa*p�[�eU�"KeX4��vskQra��[Y�e��4h���;�f��1�aDS��r˼j]c�3������8z���u��#q��CU�����$���5�)+~Wz���WG��~���4�B]�*�"6�2�#?,�3w臨�{�3��>�����(m��QpSI��g�O{&f�o�5}b&����a@4�c�A��}�V�k�h�l�iQ�UZ�)^>�d��-��.Y��z'gE��,x�7J\�R�x�r'hnU�'�B���S�h��\�ǡ#�1T[3u7 ��S�W?P�SF6�A0�*��K�r�~A4[jԫ�\�jttdv"a�))+0���h/�ʅ�Xs|�{�ؤt����=��&��_l,��[�n�T�[z~44����V�P)�μ���D V�0�����%�	����xLL�_۽ ��p�80Zl&ۃ~��Wܡ��.����x/v�	C�;��.����q�18aUB���:�j��Y��E�O6�۷X)MM��ȉ�	�9E
S#�h-�nX��O]����S��J\�\M�$s�4��[GBIipa6!6PI�i����Y�뗻���;
�4W�I���נ��,����H�A�A�_p�C7v�G0���f׭����ƍ��U���s:<-4!�
9������.yQ~1�訽y�"�yVw%�f�*�[�=��#�����ֱ^d��`Z��(�^��W��K.��8��cQ��m�SY�H�˜]V�2��V[[Unڌe�q3	��wTb'1\�e���Uj���6�b��G�Ch�]n`�,�O�/:P�[;+}]=��#�l���n}R�'/�;��0�����gy����\��I��O!j�� ��l2M�;�T��zow�Y���⦷i��o��Q����H�Ӡ�$�Ry���{}?Qߏ#16�.ŗ�1.4����4Di0��N��ȥ�7��p���}ώ���U9rpr�w��X������E�\Il"W䟀�@�iF���4��ZY��X��^s���B�)�d뺵�1��WmWѭ��-d�_��C�8����֭�sm�@1P�E�3[#1���noWoW��T��U&���oG앹YR�U[p����G��-��f���71�ja��7/'q�B z��۝�����\�̺��a�7z�㦙Q��*Z0���e�λ�����w�,�z�ݩۚ�R�Q�kE����qp�Im<ܒ����m�Y��k Ӹ�pL=J�}G�c�㙊��\T�Y��zF�X�b:Q�BcY���mA��qC��#�wێt���P���<����!f�f�u��	OA��DR:=T�[���x���x4�G3Nf�+�q�i/�r�M|V�Ar,z�#! 
J"�1d5;R���O����Πi��2��|�88P��-suԨ�q��uk�j��<���dT�0~(ـKl&Ze�9�g;1Uc����0U�]��������+Y�I1l�c�
��K�3�rH�2�r,�ҢY�	���'0J3�����L��Y2f�f&�Z���o����z����"�~Ou	�s9���^�-0Лk�Zh�IY�;V,cP.��c�l#CGu�	Xfj�.���TsAִKa�@e�����J����:��vڍ�Όp��jy�s�0fE��u�w|Z6��Ũ�^��B3G��l���_8j�l%�䏕P�w6,Fe���eL����y�Ë���c���0��Aph�h8 W�`�(@U���\�˃ք���o����t��]��b�������dt�fg����p��ڬb/TVf�S~�5��������� ���u$2��ǔN��fT��^����t�G�
6������B(���v��j�V����
���D��+<bЄC�*A�#_g޷����1R����ǜ�t�ɑ>��Uf=��ǯ6����g�ZTo���|է�>�1�x�����׹����tcqd��L���U}0UR"�ms+R [m|��h��j'ǳ�{��T�#r���ap��ڬ�0<H�ztj���;�}�w7>��Rv��o1�"�f��^��'m[;k���N��I9ݝ�ӽ�0յk�`E��
��4��>��u�Y�I�����ko����s�o�"�3e]�4��(j�3�`�F&���&�GNb%�]G~5?�]M~s���ދ˕�ݪ7�+�v/i��SB8_�LF�22Ռ���(_��	�ǻ�b�F9�u��`��釳�.�@{N���%n5���8B��5�+6M@�M�[�S]�k��4��#,u�.�^`���6=[���a6��k���A��=�B��Ԓ&s�+M<���3���&��}�&&�Y� U�Zci�L�t!&&���a������	g���o�#"I�5��D{�By��t�R;�܆p��,�������Y��ģx���6[����.x��z��s&����|U�nW�ٵ=�޳=�d�j��_[��Ȭ^��v�<��r�<*������j5b��z*��A��p6��+��'��=�rZ��*np-6�K.�ɔ�s�y*��F�Н��p�lk܃#h�%�Y=��#�ߏYb�f,�m�����=B�)!�k�;Ƀ5��5���о�Χ��S��ȡ���k}��#�c�+c�A�P���5�ve�#l�ف�|0B�My).3�8.R�}����}{���>�����]���윓�F�����w��u��GF�r�v=��)���5���X�ʑ#��Q����:�*q��7в
�ʴ�o�A�)�`��?Ĵ��v������]$��V�A��8*n ��m�m����'�WwM�曩�����w�}����R�� ��5���F�_B���ҡZBL��*�\.�Z+��QU�j�nς�Kw�S�>�}�A컿	�l͖��B�^fI1E��z/϶
����b����1s\��Z�{��;�,ûS�{��l�ʒ��93�FpɮT�s�Mpǧ�.���f��n	�V<�f��u)S3%Mڳ��Ô�`���F�|3�ӏ4�pj���w�b�P��y�a�4t=!;�<���[^Ӹӓ�Vc��wQF�T��u ��E#Ɉ���#K��{\f@�!ij�Y�f�jl6�e����;Y\k����K��l�/<]��
�X�jһi)pWV����v��8F��-%L0�R�vf�6Rh��!3#-��ڴ�:k�iE����av�[�4�:(�E�$%�ۋH��& �e�++��a��n�@�Rk�D"Ytכojl
�iJ�0"�Xa�(Z�ǩ5�
,ؑ�r��Y���u;UV����;�2h��m�c�FЙ�-��]��!J��r��qp���6�����>�z�7,ɩGa�hV�i���0�U�-�R�[J�Z�p�&�u�!��6���4�aƱ�V�~����֞_js�7�/c?2����)�K͓T����:J��Q�YV��gg��7q�ٳ��X�;&E#{��`z��K�D�-E����^���@�I�/�\]�"��Z*�T�2��jg��G	AWɸe�����W���f�v���YU�_�q!B*�]xh$j��ʴZ�ξ��$x�R�BiF�;����f^��T�7E^z���u��Q�}HCt*6Kk�Ըҵ�*w��#�T>R�CWoGH�T��t�P�`�@�I��$�nG�*���Yk)�r��̊K

��&�Q`��Z�`��]��C[⯳��[z�>��  ��W%�^GWM�~>�8����nV�
4�MQ��{x��>�F�K9�|���ٽ�ƕ
�U���1��YH�y�p�E�tDߟ#
-M+������������eZ��-Y*+pA�\�ü>�w�Y�@xT�������EGmv�er^-ڽ̷�'obQ�����w�b�G�}>��(��X�ҕ2[���?p�՗l�K�d���=~]�����l�D����.e���JQ��ޏy�m��ZVe��ndFY������C$+D
�\&���6��&�~j�m���+�/2j�r�4�yL�X�ە[y�!k�)�C-��b����\�����k���-�r��5!)t�4X3h�su�6<��E��Z\�<�4�-�2Ř���߿ϵo�U���=�WZL���ش�H���x����E/a[Z_�nDV��[*S���]��=д��h���gG(י���p���|��^�T���T��CA�$���ChU���]	��:��5�����{��Nޕ��F�_����bۇ�"ˊ��iX�r�q;c��v��q[�ޗ�
.y�^�r~��Ԓl\8��R�H�N�h�(�B�-uw��M��"�����ꚁ��Dz:EBH�	M��N=~W��#Rg&i9��<O��-�����k��/f$S����gC[jj��J$�}���$���K��s�
d\�䉋9����ؽ{��U��o���U��NT��;�äBJJ��~z���<�mc!p2��w�~t���b���QAW�4��� ���t���,}�M��r^�Op��J��t]���we>G��[�5=�����%���q����_.��L�"�a�j�r��R{����hu��5,���#"�z���5[ �i"�%	����yC�Q3"�]h�jf�)\���#{O�#^v���F�FH��`�OR Y���s�z��|�떚�c{qX54^EH����'�=ȫ��U啞.p����F�k��k¤�qʄ5���[��������L��,� ��\�hұ�l�*�Giz�ۅ1J�b�Ԁ���f�H.����h�:�@-�(�7Zf&cfp��s�@#���G��+^Y��V��Cʛ8(�(�Av C�&��;�= ��v�[�П|B5_��1;K{ ���j1��y/t�v\�R�'�4�l����-�*2Qay��4�ȍ�L���6��<9w����yNb��н�5}���̿���O�}Ҧ�]8��e��{(�wڳF\[P��J�\��Od%]���{�QC�V�׷���t2�FI��"	Nnj͛Y�f'az<E���z�7�mlzc�
���>���p7�����ja^�վy�F�����aŻ���6%��p<�ȲlDN�x��R��*�lƐ+w���u��o��]��΍��C�Z&��b�"q�����Q��Jf����#�3;H�P9G�AT
�
#�����MЬ*lu�O/�<1粧U����y׀VkE�%�;���sk�̰h^r�h����a���c��F�=�iש��	������4ͽV�闔_���}݅g_X��w�a�Y�@�S�<@���,=OY��C�$�"������A��F�ʁ�N&�xʋ8�W\����szM?}^Q��s����ul������WOk���}�r��mfR�仵v�V�:�Rs=��=^�	��2��e��L���72�#���D,����b��G56�f�s��^ll���Ro2٤¤]˞f(-��n��Nۯ{=��m�s���&�T�{X�b2uV9��E�9ս�~�_P�ӺǾ�p��Lvm��\����n� T&�)Z��,��㗙IayQ�>#1�o:ͥ�Y��'�-��q�5c�)j�;����۹���(S��X��8<�w��2?e�IYp��y�^�)��o��,�/�Q��Xk#���n��>�<�W�s�'�}�30�ñr��rp�kq��U��e]{K̵ܐ�+v6J͊�pdn(��7NV��̸Z�nb��_|���|��BM}z"���%Qz8�Nةɒ(�w��碽檲t���1Z�ԝ�������'9~�'y���q�P���X����~�9GL7�4ȹ��� Q�	(��e@I�a�}�٬\ݙ^�Fr��F�y�L�>������βѼ���i���o*�}�[B�������옡ݺ�n�{�y��=�y��>Q�-����݄����|b��˒�Aك1hf�H����H�����"pB��j����hh4"����Y2�QQx�<�ڻ_F7ƨ���:w�뾭0��V"r=�E"�d��^s�a�R�f�B�^�uq���� em���wd郲��n�̟����e#0��tn��3;{���9��������K����诺}���fT�i�k{y��s֧!���n4�Gv�{9'�o����y�wc;Ӥ�U�p���:��6�#2��{[�!a�9�����:�8��������m���p��6Y*h���mC��H����r!�g�
vr�:�a'h����@��NXK����B����=K�C|���g��힡b`V�������*a��.%���m��Ҹ�z��8�-����Vx��lU�\��`�-	�)�\ӌ��m�-�[��J6�as�mB+k��f[E�].Ř�͕9�6Rni�E4���n�eP�Xz�{�k̗uWu�H�m19�ٺ3"ڒ�˝}��d^�aT��x*���Tm�pԫ�}5�HϪ�K7�KמV+�3���-Y��~䟐ڒ�W�k�����r�@���ۻ>������{�ZXi蠅3't݀�s)˻��5n�e���5���&k_T�m�=�_p��Pk�$�Fwr�{�n��h�'���,`���U^ƕ��>���w��1���A���)Q��Q	��P�-&�IfY����c/~�>���q������̵*���mwc����}̢D�@Z��Q��?��K�Qi��*�+�2*�W)��F��/�/xp��8	��H	��vn�)�VNR����<���c�&=��][��K����O���y�8^h���2���օ��+/;��r�����AZ+M"��]L#熩�F�����vl�lm]L@����w���ǣ�Y �\�6��	8@��bݰ���ea�+E����mfś�}�;O|�}���8�^�(��V�9ʷG�Y��4�W���LW�D��H2|�8�Q��x��j�"陶�@܉A-5�s���nBѠ��u��흦rx�iL%�#��u�j��ަd�TNSI�ȅ���NFkS��1i��)A؞�O���߫�ᷦf�ˣz78���� �cPxlJgiڑ�$�&vr�F���w���b��q�{NLɎ����[�)
R��i\=�ۄ�/^�/�<�p�3c/�־������Jk��ë�d�\�hp7�����nڕu�X��V���k�Q�fSaI�h�]�ږ(n�nɨ�E��v��W�$t-�m
�ܺ�-f�Ws��3u���d�L�p\��(��4 �d�������K���\�-��1.�`�q5�wT!5e�n�����U���:c3;-&#)�±�ƓJ]٤̊ ��l��ivB՚�(�⚺� msqi)� ��f&����D��i5�������Z	�qB45(�a��I�y�<�x�n��=F�2�heY������h���E�Mֵcx�W��q��օ�$�R ���Ha�i ��u����� ~[}�;cW8���FN(�숬u��9����U���ᾨumM���{tq纕��`����ǶS�P�y���oz��d2�
D$_���M��أ�UoA�(���@uPOk�<�]M䡷�I��Vuj����Bz�W��s{� �I;���H�M�k���'�cW���A+�y۹��+�-�*�5󃫝'>y'3^�SG���`6L0�2����1E��#y\�OX��+�|=�1aw{��;A	�������m˱������]z;-C�y��s�V
[*�[PkJ�cS�v+#��=�"�ٿ!o`A`	Z@&�)����U3�{lz7Y��pj�}�&�.�6����ڹ�~gn	�Cס�5��Ny��W�-�n����q�[ -u��Xnƥ{�Cﶻt�EG���x�O#���~��֩Z`�q��g�S�}��[��{�/s.r���®p^ۄ=����C�����&re!e���kѽ�1R��@�0Q<UƉ~�h�>���ξ�yCe�s�D�86c�Ȩ�n��{0��Ԃ�d�Jc�?�mD�Rd��hY�*�m�e���M�fyԉ��C�S\���n͆�b��QM Ѧj��!����&���a�q��dh�Nn��v7>��%q��\��VcXL�T��!��p�ӽ�S��U�F4l�T)�hճ��n�WG"CH� (a��jՕ�O�M�sx��>���n�+.�B���r^�v�k�ŉ�k�oH�>�qe�G
���ޭQ�|7�s��n��wO�-Y���s���i�)��^G�o�2�Z(zF������DG.	��pHp
p�B��;�s�<v=cو 2�V+�aX}�r�K�eh�6�Υ�yϏ�þ
�πǗr%�7�!vؘk4v�fk����́���Q�s���U��GV p4p�!�	�6R����5�s�f��?f������D6�V��cZ�]����R�߅�373���iïy�蝓+�c��%�p#���.��`�[ �{\���)��<$g���{
!�Ii��l�-��tT�Q��ͺ]��3����q�n9�k/@��&�.���!J�=c��%���8!L:A�|WT�f�:�g�H�ص�H��ҋ��r�D]�g��Z�D&�1�p�ٰ`�ͭ�m�F��Lnh�%]j�b��4�˳����ъlm�WFm�˂Sl���txPG8/0W�-[��#����d���s�v���̭7ZA�CGۑz���� }b�4����9�D�	����X����S�:��)�Z
��J��L�A�	�f89�3'`��<6s��Zk7d����a��.���Y�tf}6�X�����Tܸ#��]�_c�1�P��gx�݇���0���ϣ{x8	"�d�9�M�yO�╳�(
�4�.&�����z�ۚV�fi��̬�j����>�T�Kg��]Y�M��g�Wʝ��!`�yգ�ӗ:7����3�2�+��s�ҲjP<���/̈́�C��ky�=�&e�!�p��a��%;�KY�ɥP�]�-9�-�#hkⶮs.M�.<.��U�uf�c��JY2�_Ԯ������ۖ;�nd����T:�����i��꫕&r��|���Y�3a价�͹Q�<Y[T(Hs1���N`�i�ɨ��k}�}�H�s<D�e5i��`�ej��2p��RO�����[t���W��-�spL(m�d(C���y4s2�ى�^�f�<s�v�}���jD�Mvz]_���h�2�؁�+�5�ӄ���	���u}~g>۾ݎ���^�w��T�kf�K�=$	}���_�o��\���Ľ�T�����0<��A�Ai��rwjz��h(wBd�+�<Aky{�
s9�\���"\�P��|w���4w��]�Oz��=�,�u�����_��+�n����p��vg�e*�t���V������F���]],�6!�fF��A��
3[�f��z�3f���]ִ�3V����7��s��|��e��w^&%Uq���T�$c�7p�I9��0�fu��߻8I3��^�s]�2���O������v�zU3#�zRWJgy�	��JH8e8)��Y�'A�^>�E��4�4;�l�<�0Vq��5O�z�P>���}���yf���r�����u���E���|\~�}^��=��vI��kQ�wI«��+�v=�ُm���v�Ci�a����,1��s�
��T��W�ލ9�ަLO�w�Ȉ�g��Q-�V�iG�p.�.��S�Iľ �t���F���0��'��r��dI&܊,��"r�˓��у�o,���Cbl�x�NE����d�9���ڔ+qd�V�������i>�ume�]t9Zb���K2��V����v�ν�P��E�rB^��$��y՛{(�|u�,2�t�5m��{�7훍��\a��l�� "��J��d����+.f����݌\9 r�*>�/tU��SYWtsp�u�F�q��T\N��7�����w���C����E<�˻�;�}�|U�2_\��^	����o��+�3hܬ���EJ`Ub���抲�l֒�`�L[���b�c�vv��ܳY����4v��EJ�هbI�����ӧvqh`���fsnN؋��w����]j��Vw�+29���]L]Vh]60Ŀ5|�=q�5۷�ӿl5$m�i�j�Km�&A�*&fD��U���m(�Sp2��d`��-B�<��ۖ�|Z����-�5��h�_f�9����f^OVG@r�rH�r�g	���G�wn�l}�f+JO��v'a=��5Ĳͯ���W���Ҏyp̾�z�����$�_F�_�1�.�+�5���ٍU�����8<����<�hz͙���S�]��T�N�3�݆٢�k�(�i�K���T��^�Fq����-7��#j=@X%�N	(��P�
�T�3��޸am!�w�.K�X��.��^��9�\�E����>!� ���\�5�5���\j�g�5����ռ�K�vQ9+����v�y�#���݇����$t>���E�Yi0�@��Pl���Wd��?f!} ��t���{Rg�k0Ez1�5�ev�I��>�����Lr$���dT�]Ʒ��M2;�����-�Qc�;���?��'�^X����}ɥO�&�4 �6k�T���\��i�ݶC7���;��z����7c��&�aO�j��Ԯ��]wbe'�F��h5ަf�f�4-�����V���Vd�d��Jt���z��?`xGPgN����cWk�Y����Y�T�Qۻ�e�D��,@�jۼ����v��O&�$�ES]���Ӎ~O~����-�.�-������v��]�Y��W��� SF�l���Y�ԁ���v�؍	����XZ�n	�&��㭀IXB�V7BսIq��зVe �e��jLQ\^Ɣ��K�a��B`&�6�*]Վ%ֳlM6�	X�F�&J�-�$
��h���񲐔lh�X�՜$k0�s�m*[2��㵇T�6K�\2b�6�	S��m4Iv�sa����S��-�A��G�_]6J+��(�-��9)]K-��9��m�nW�����t���e��˕�ؗ[Flj޷Wmn�nuh�6���f��z�i����Lj&�m��錚8���n����Eh�����l�V�ʉ��h�!�����������;�XұG2��S�o>N�I���͸����z|ໆA�>I�w�ki��>��˶ր���
�2��0�I��O�2e2�ٛ�ҏ�"�o{b�R���_,j�ؕ��+�J1���m�fo뿓����n�����)���f^���=ٰ`�з�FG�2�l���/�*����4��r�뻻������]��i�l(e��6�_k��z�yc���Ϫ/�|+=�;|{2.sjJ(^f���g�'|\��fUcEt.a�=����U����=&��������z��!zI:�,�	��0�*�M(C�|�^�&�m��᰷hwt��U{��^�uU�}&0Ol�nײ��%FX�׏��y����=�*}+M��f�FQ�~	�\p�-�*C�Vz�U� \������qQ�UYP/�_�\����T&��H��h�/ ���9�@C����4����)�zm�Ca�K��-��n�·H��c;}��6c��5֮3��=�v#�z�a�{����x-H�*b�M͏e�|jr��Y }P "`��� ��ř�rb)��e/lk��,Mf��l�L7\�Ќ6յ��ca�8J�ƕ@���RhG&����Wx'�����u��>�L��^�jH����{��n�]v�2ҙϝ���[4��M
?���ڟ8A�e,́"a�k��$�!�l�xı1�f�oӱ{TqH��=&%>9��5�8o(�/T,yE�~�w�}��+��9�����s
���Q��p�:��ULS��:}�^�]����A��o�P��a���8�gtƞ�]Ə���!�a�P�)�G7�;����Wd,�����N�==���f�w�4���Bĺv4y+���9W{  ��o�f�&��e4�{��K�F?6��ne����V�'J��!k_|�w�YޒK�|�ʙ���11���~0�_��[s��r�ϴ��pV^Z+� ��ep3��
���DFjS��+e����o�������S0+�țƲ���iw�o��y��鬞f��x�$A���B1�/��������>���>~��F]���W�&?��o�б�;��ܜ�ͧ,���Kp�������e��a5'6��x��!m󞁗��N6x:#e��^t�����`���J2�J�L-ՠ+ծU��K-u+��9;H�b-ѭ]t-"�4w8���&���	�[�pu��n��6�Bw���>�x���H;
���6^�[�5�ee����n{�o?hU���Wo&]ϼ�6o.���j���e��b}���R>�(+��PR]�L��zO�����߱�'��3�~ѽڧ�v:R�n��unlEX���oZŚѬ��m�y�>�ݴ���eq��=82mh�>[HӠZ�8�-��^P��&�_P{7�c6#��wUue�QV�7�*A��	Y�9�m�0����{��0��<�9~Y��K`�yl#FFkʮF{RK�qܯx�Q	��Z�X92�`���՗��h�껮[�\���Rˍ�#e�G[۸s3&y	�1�+-B��.��)�1l�.�d��_�T˺�@���>���:c[�O�[P�R���bډ`%��Y�F�}�^�,>zv��R[���r�r�4�����[��Bl/����Di�)�yN^3�{�s�fe}����2N��ޛ�w��,-Mg��ҢN˩��=n��̥/�7�c�!+�yG��W�X$&M�Q��v��<q��Mn[bҧ�D��Κ�;5ѻz0�v�e�DF�^�����ݲ�',��|�5��T]�y�9u�MJɣ|}Ks�97��k��ٱ7oϮUE%�mJ��%�T7
�t(�[���}~����$�]�u�7ԗ��K��EsJ�qX���wRrvd2ԋ�`nn����2@���S:�`��ɝ�Z�˲f`�� Q�^eD�1����E��,��l9�7sK�k�V�9����33��K3J8QtKZ��j������[��nܘe@M�g�3����%���R�qd9����=:Z9"��a�w+mv��M���a�y�������j�ݾX˾�w~1sP}�Y<T�8
��,�#&���=��[��U|��Ϧ/Z�:ֹ9�SB���E����7row��qɩ���1�^s�mdb����k�Ѷ{�o�^�fS|�_#_{h��0'qIo���ϧ��½�Jt(l��Z	�a3��}����xU�ֱl{+<,�wvtz�OUe�^.��~�B�5tE����,���$�m� 0Is��{�}q{:�T����vR����8GOt��|���IuUK����wǓa�h	��I�_U������W�.�ok�V#.����$��W�f�w�n��u������y�$y#ʝ_�I�TY�1M��w1u�=��ɜY��^([�TB�y��q��a�-@M&�-5\����G�IF�aǭ�R}u��<[�jy�V5�,���TfN�tW3S'p�QG�U �]��s�{�k�<0\�T�o(eA��Ø��Wgb&�f�}y����ܰf��1�&��3Y]�]5P�f�k��J!�WU�n�Z�qv���e6�4��.�/L&�-vJ!�U:�����X����D�g�D��+m���96�7g�Έ�7n}FG�y��	�������{7P����{��L��\��ȫn�2�nC�[%�~��0�hd#��'�Gz`�����7����k9��^@�D�c�'ks�<i�����vW��l;�W9��l�������L�I�7��ME�W^Kw~�ю���!^Y�� x����%��p�0�d*��:n��M��re�\��D�*]mO�Zg��6^'j�N��O:cb3�����/+-d.��J��W֎�h��jw.[C��6�W�c���J5k�����TRP�eC.���������b�H�m�*�������Qu��Э��X���Ϸt��Z����T��g#z'�)���Į-�ž��e�B&k��? 'h8 ��%��(!�YbO,�����Sd�tE��=��=�ng�������,���N�h�Ε�e�Šu,���6cfn�}�T��7�Y`=�W�9f>�c��:o>הYC7~.-S�J��|���ׇ����PE�������N�Q~OK�p
�/?��zUu�p� ���m�y�C��v܀CH��!8x� �Q� hB�(B�`I"+&T�2�L�HJ0�v�
�I&�	&�OIH@ 
�H� �HHl�?�!���d��7�%��N������H �!$"��d��*�e����-�����庰�mq�t�*����}�����QPqYPk;}�?;����I]�+���`Pv݇A��I�I,W�5��-������=�x@UE���k �
����]�:c��!����Y���#�A��AO ���W��=0�d0$ڒ���:���o�U@�-��(��n���VV׎6�;�l�
P���A���O�4�?����M���QO0�N�f֩�NeN	�c�sE҄��4��c��4J���^9��)Q�
��z	Z����e�3��N��ݏ(%�h
T[�u��P�D�5���mwM���AI� ��y��6���`�w����q$��±Û����e9
��~4�)m�b��&���9t�1��9�^!#�RM��e������R��]F�����L&���Jtg5��W��y�;�<��ڟ���u��~� I,��� m��!�!HB��$�HO� ��D� @"@�!� � �$�zk���|@̹���a`\���b`Qt�"�*$��΍l�cz	5�N��2	���iP����K��!�$�
�v0c�DAjw:vK�O%~����V�=!�Uk+����ϧw)`nhzƇ8�w �1ߌ�|���1PEq��#�Lz�H��A<r-y�����}�К�\*(+��W���3�쇞f)AΠ�/4��PN�@ $��_�1?���~�?`�>d	I@������=~�a'��C�`7�,�Q�h��<58��ѩ�	�P��"+)XAq���~ŚX ��D��+G��v�����}������}��
#�l��@�?.p�0�a)����K�o�AfE�!	����+���oǼ��Ky��@q�8X�\PM!��X``�h���/��p܄�8�p�q�[�K�-x�m+
���P ���"F��0̊�&\�LCD�HHs�cͯI��@�{��P��\V�#jx��]�*���!��.!����Qv���&�풕�5��E���ɶ�+O�F�D١�I`WF)w���ܑN$�� 