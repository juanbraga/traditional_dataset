BZh91AY&SYX�9a Z_�Py����߰����`�{�"� uWz�	�� �i0M=MF���F�44�G�L���h��RR��� h@  UO��T)@  �   )�$�	1��&j4hш4h��L�1�2`� 4a�S3��������C�ɦ�<��I aҁV�$� P$ �_$� $�p{�����$��H<� 2�?ٸ�bH�Q���dܚ
���g>��rᶖ��%
�  (H	PV�����   �	PM�:���Gߊ�F�Lw���j[�T�'S}K��Z�)em�F-�`��bS�r����"KP���(&	��9�"!���|�0��<!��\���[��:oR%����Y*��++zXJ1BC�#�DD?! ��R8�����M�_n-�g��KI$�X�BI)I'I$�$RI%i$�"�JIJI(I%)$�A$�J�)$����������� �q��<�	nT�]�j�N@/K_6�OD���FE��b4[��I$�B	h��+z��coJIݡ���c,:��M���{l�w9�s�<�b8�9���I'�������C9�!6Kc��+b^�c�� ̐6���\V�n Sei��z�:�I$��f�iq��yЂ����[]�-�e�:W��c�6��؜1ۀo��s�#�Y�I$���Ƴ[��赐&Ƕp*ؓ1 J�bx:d�B�wweI�-�7:� X�C��e�I&�O�)�~݈$�9��p,6U��� ٴ��q�"Cp2x�n
�(�:ZnRīTܵ���Z�	$�KN&43lM���ؘ�ё&��w8��j4=���U��w�TU�əm`�\�$�I.�U����Ee����6���/���R�`�.����J�S�¬1�b�k[ ik�/v5d_5]zKl���	������lևt��1v��w%� Ʃ�jm���'9�s�ٶ)�_l�1�m�vǹ2�[�1L�U�l��� ��o4͕��3�ı���QlVk5���+����֭Ų3�O/c���G���ަ6�� �d�w�	p�Zn�R����Y7��V���D�AB
 ����(,�L ��(((("�I$("

�APPmi%���9�")�̐A.�IQ��d:_0�*�;L}���$cg2�`�{��rt�FR�N�hy������|���"i�O/&�r�2l�q��N[�6݆���Q�̢�R�@�L��#J�4�=��]+�ׯ���s?`�r� c/�\c8bQ]|FQQ. �WL��ON���%�� �VZ���`�,$"��w*��p�5����%.5��"�(��0����g�+)o��-g�{��h�l�H�(��1ZA��T�E�|D	��!���Ϩ,
��� �٢9�<���UB��;K��m�����"�:t�� �&fW&�du8�59��I�R�5M��D9��TL�酤Q[gFU��cZLD �z���m6����1R#��MV��BI�.ôXB[,='�L�\�2z�$-��*d
"�J�Rh�K�!hd҂��)����N��.���,ɑ�����1����!���w�}9�3����`l�2%/�x�y��㸷 @r�W-caֲ��o>��1XM�`h�1@�8ƅ�6@ ]\+S�ׅ����b��1dE�d�*��g �a\�r�m�1u��
�%F���(�&_7L*m��[Qb�LX: �;̲)9I�L�p���^��b�K#}rW�4ʧ�©��P�E4O�Z���:��j�`�VxF3�<�f��iT��SE祠�h5��%����)����