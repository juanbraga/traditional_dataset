BZh91AY&SY>�q _�py����߰����`�u�_x{�G͠m���H��<�����ҚyO)�� ш�114�S�	�SD� �` =@0 OM)��S�4�6�@1 i�@  4Њj=A��42h�ɦ��$�H�jh�z��茚h4 @���Bi2h�OI���C�<F�� �=F{��CH��l�H��ns�RI, �D����?�S����y�#�~�\�T�#�@�,�Ҽ�����s~FH�EU0�FUP	Id$�*�u7�%A��	�Ð)�B�
Gj��&��$�}ǀ�c��N��(�<	R�I%�.
HQ�Q�+;�v<R1X���7�22(L�Yh������P5�X����Һc��aH�h �H���/�{ �a����	`�`{j��wJL�	�!�]G�Ӵ�_(�osh��(�9B��ڭsa��V�V@�R�R�ր�mئ��a�
*Dh�c�^;d5��
]���dU-�灪:�ָ�4�hE�A���wG�B,x6��.�V�:�Fw<:�B�k��ֈ4z�Z�k���&�Lm�����*��0�r��\?m�1i��=N&�`[�"�n�-�Ô�QIw��4`��c-,�IRO��N�X�l;e�k2k-2���Rh��d�~o`�G@�THB����d)UF�`PAS�rK33�YNܢp�2���̯34L�4Ӈ����C�F*��a��bh^mHa�F��˕�jY/�B����x�l�¶�;d�0k�nޘ�-��0yN�T;E�ec9ܾ�J�3�/է2����GS:�m?y��K�K5 ��X��f5-p����gjq�._%�mV�����2BBH&� ��"�=�jO�'	��(N�	.ĕ����T�����!%k�I	�a-dN�%XrP9�KPohQRKZ��X�Em`�nU�V�[���M�����8g��G�x�Fs�0,.t�T��H:�t�����-aw0���쬙����Ȍ藡#�G
�I�� �ӛ��R����m�6�dΟ��U�������>Z`��'T��S��y��Ai�����Vp�L�RX��)�:� �~%7'��>]�����vB^i�-�6��`	B�ꧯ�0��+� ��e~kp�����νJW�q:I9u��{i/$�� �� P�BKO��\H��SzLJ'�V $��څ�A*��%x�{�dQ�����P��ԑ��.�z`[A�ȃ{�ŖTK;�6˼��]Mbe�لmL	'��A���w&G1��N���Dd�u�-���6�2a��Q��\@w�D`h�g�s��J�4"����FA:���b�Uq�,(�P��]��N�d�r. ����*��E̅�Ku5����28�WJ0��	�SHjw�*���	�қ�#���6�i`�N�����j��l��I�6*HR��g')n� ���v�Z�Dۗ2� �INs����D>�Vu/�L�{�M(mRf� �9�f���V�gE�h>�S)���z���nra,ɾ�L��fz�(��,.�D���&����&)� �Z�y��>��_�M5꼸a:(���Hû�"ԍc	X��W�5z
�5�}m��]-�*X��~C���0z����rE8P�>�q