BZh91AY&SY�0�� 0_�Px����߰����P��`�ܛ�.n`�H��i���Dh�4hh1� h%�##J{Tf�zC@ h  4	���Bz�S��B4h� ���& �4d40	�10�I�f����F��    �L�U�����$��K��C��f��d5�~h�5�#�Y�������X>,�l�4�+�1�
����q^FR;r���m�g)Di���y�H3,ƌ��)�`��ؼ�k؈�R�Nݑ~�1<UTTU�Ƹ�A���T��?��dKT@=�HѺ0��v���6��0Di�^�Y����d_'�1�F�������������m�p2z�N����b�8-I�(��o{��f͌��ĕ�8��0/(C�1�
���y��0�}��X�鎇~b�B�e�1��yf��}���=�h����"$�~-��ߦ���H�ؙ��ٽ���X�F��H����R�U\�*�g5�ȍ���8f��0�&1�x�'D)A�:E���B�+�bq/��N���1�Y��� �qs�18kz�ٺ�>~PXQ��&7�lyp�3x��N3���<���i�BC'8�j�b�6EI��c$�a��0ļ�:��['%��IB�U0�,�q�a����-k�=V��j*�wVG�qF���#�Rp]�&)\�]��I��^�Y�� Z����+4��F�M���ZT8(1�*����0�rY�u�d��l`Ҫ�b�%���Q=�jJZ���)2�� ��3��T"��T��&�	�KV, ��X��!�WIz��a�P)6_6��n����Ia@)x�m^�%c0bPR�9�F\����j�Ѷ%�����l��*�[�DM����\j��Ȉ#N�b�
�R�S�A�wqҰf9���p~��I�e�*B�i\Vw"�E¥��ER`���HF��-������P���,?�I"ʘ����s�,<sn�J�U9��r�~�2�^O���Sd�d�24��r����)�	��H