BZh91AY&SYM�I� Q߀Px����߰����P>r������5S��2�F��I�������& 2zC&��L��j��M��d     )�)���������Q���@ ��=M=CC�0L@0	�h�h`ba"S ʚd�<��Hz#L�� ����E�H�E�P$���z�X�kv�!���'�!*�6�FI��Q5V��/��i�ɹ��F���r}Ը�h�b.��s�?�5��%�����ӵ��	5��a.P*��@��yl@�#�����~�k^�d����g7�+r3n�2���:\��D��;��ͤM����@�W��s:bQ�$\ɴ5Hk�&Q�<�_TԜ�֕�)�m�[���ߟ�hI		+�Ia8����4�:$P�8�yE%�F���֏( tDA��ԭ"�r�1�Mp'S�� �
&���65Ҍ&�����|	�}�Yд�m��d/�Y��t�_�}DIecU×Ն1�LuӢ��2V��x���p�Q�\O;ά�2y��ʋŽ_��8��q�?XB(f�0��s
c!���R�%�3�mp@]D3`��/�t�ō�n"R���p!�l�3	�2�:�����@3�M���t�^,�H���Ʈ�"Fe�@��8P�����Q
�h���8�h	�9��*�e��ѐc�/-�Vt4^.R���Ww8�6�Sޜ�U&��%̤���y��`��Dnˤ��`Id�&i��P7LS���v#8�p6�<�GvU2#�ɓ�\�SU�$�9�y�	j�ٶƤ'��9X��)c	"��� ��;v��+�q�;#���$�04�O2��3�G��m��v�,;�WnJL��	�J,��0�D(�@����膿M(9�����#@�A����b�L��f&%�0�r�Z9��2���]B1ԣ4A�U�ñ[�|⇧3ɜ���_�%y�qT���^{��2,�B�Mߨ)T@�� {�
v�D�8"Ņ*3�u��]\d��8�ȫ%( tb���
l[���mT�܊���c�p3/�ħw^m�8�i��_�:�ܑN$aR~�