BZh91AY&SYb��� 8߀Px����߰����P�s���L�qUJ"W@I�I��)�OT��FmP�4h��4�51�d��G��Q�L��FzDL�G�h     4�	���dɓ#	�i�F& �""iM��Q�<��&2zOPz� 4h� ��H��Љ�B ,�(B}F���7U�f$u�&��Y����$���D�	\���.��~�.�w���Je�nJ���t����^��rɴ>��Ev#+%U��a��7-2�󫹬%�85_��)o㔥��?��jP�Q�(a1O8���D$��i���a�( q���><j3&��5щ�v���>ʒŐӫNgW�\%�r�������le`��Y�.D��ewJ,Beд�R-���K%���#k�4��y�ɚj�d��D�lYDV��aiJ:���K�X�,���N��xi���tШкqw�Ôe���1��n�/s�Ƨ@v�70�gW��嗹�����
�g}�̰c��-R�����6f;����eNy#w�tŮ�r˗�}-6Ocai��U˭���A]���st�i�Lg�����:�8��������`�
'����2X��ܼ�U-V\Mv�N��xo:i�EĒ���%�M�� gKEj"�lY"�e��d���5{Uسk @�f��t����/�,]�}�3�����%�(�:���|ۗڨ ݇��F�G��{�/���?���Í���v���K�����L�D�y��Ӫ|���l5���R�]�a�K�������i+�V
�6 ����=b�r�jβ�J��(��"�9m_A�u���xn Ur7#�|L�[���^�+n\A#D���w�І��)즋a5�Ve�x?E�fM����̓� iK�0�d��[�Ss�Jh�L���!�&N$
5ܘ�(�*�J�@�Y>*��*�����G�߰^nK-�� �(Z��V�
oF��ѾƳԎi�4�V�,����qY��++�K_0�����W���̘l*ho?�`t��}P���6��/uy���m \�p�tf�
Wߩ�"�.?s	f(+�NQ�4@��J��JCR�_R@�*�7�� ό"���[�U�U]%����K;��1p�B*/8^i�1�ƒ�d ��%��I#@ip���u��}k�:Te�� ����O�p��&A���p�])ZX�ӋX�p��θ� ���
g��e�3�e�dXu*b�H}����
b>�Kmǈ:�����o�B��D�I�To�($WcDPL��l�ZZ�Xp���R��l�vS�Y��ẅV�GT�^Z���[���z��-*kK�;Mx����2R�����A����ɐm�۵i?�w$S�	)+JP