BZh91AY&SY�2�� �~߀py����߰����`q�>�r�I�T�R�IA}�      0 ���A���]�rk[P(�*�]ܬ�j�;m�˻9� �JJ� t㠑!bJ%�bJ��mJ�TQ�d(��g 2E(+,��(�*Qf��(�%IJtҸ -)T�Yd���D�%�RH
�)$�D� @4(�h�35D�IډJS Q;�O�-�h0��E?U)I�S�A�� �  O�b%UMS�`a&&!� �MOS�M��4h� �4�@S�j�U20 L      �D�4�M�*~�I�OI➣FQ�=#�@�II�i'�������  ��pjs�r�J1 R���ʠ���h *AE3�D E*!(|��G�k�����H�r���)�����΀d=��,�ﰩTK��ݝ{s+�����[���Y
�LaLI��T��+ (���BVa��I� b�1��Āi��B�Ti
�1!1�bI�cHd�!
�d��!XH�&$���@P���$P X@�AHJ�!P�B�� i�4�Ad@� ��,����Hd XH,�$$��Rk\��S�,���?���a��>�O�g������~O������ǜ東.$	� Q?F>��H�e �JT�VkK�f*�L4�Q7�*sV��h�^'�R(�xQ�)Ea5Phȓ�Rˋ��n�d\�X�aN�K',B��H�e�L%��9`��T34�}�d7��)<���EL� 9^k�3��+Y4*%][�!]�A������
�F�E՟���PMH��QGl��]�*��/t]����6�&�����)�q7v�6,E9��v �BQX��AE}m�7dR���!��$ܩx�۫M	H;�!RI8%V*iMb�*�!�%	��&$���LY8� YXY������dʺ&�pm��$ٜpn�q0d�4[�R�t���jNdb�&2ʩ�S���g�	������y媺�Q!�n�����Qg��X�]SLB.ʩYm]9��KJ�D�!
b��&S�7W$���Z�7�����l�S9�\�V�$���a�`Ŭ1҉Y	��@�n�X�R�+B�8�Am�Y�LLLˉtnMJ��.�)Ta�P��!L�qJBl����.�(.�*�������0̕ݫE^Fѥ���锫)U��`�4ջr�3���V_�

˷xŻaD���6�� c��&�0���D+ȑudĵTfX�u�e�j`��)�S�M��ff.(���dH�`6i��$��YF�J��*� ٻ�-�6f���2̻�n(�Hd3nDY�DŘ�b�t�5B���,EѕX	��8�ɇX�B2jT<X��P���FU^e����'7����!�˒hed]�����$�72��ؗń�\T��UK��E��B��0��bbԔ��LD�!尰�d��ɒ�s8h*x�qn�)Pe�'m��e�h�k%"��72�G.*�q5bJb��`9�7m����Nd�qf�H�ɹ.�đ8����ZF�Ƞ6lX5M��G>�pe�E��8X�"˚dXs�.���C���eڰLa�J��UX���*c) 7J�Vd:��8�5-a I��dB�rD)���s�jJ�7r�Q&*�m�B)buZ����\ؼu)�lD��GJM�S����7b2,2R��bq�T�+WxC�LX�O)�ZS�X�O�q*�3�(�ui|3*S6T͂*�%M�ByN��7��TW�˂�ȗ�Fo$Dc��P�b��3@�B&de3�	6\ZVқ̉��k:����`����� 
V�)�C%�MD��U(O��2�)��у.٬H�C���&�
T�ī�2I���vרuFY�����׮��"Bݻ���X�C�>������7��p����������t��{���f.�g�Ѭ �]�њb]�I�c<�i[-��ȳ[��ܙ��4�5����ƅ��X]+��\�贏4n��Ggj�m�F�lB�FT�@,V���Ƙ&j�)s�n4�%�і��D�
�h���&R�pr�MMF�R�l�F՗-,��s�n��SJ�$!��433�)`�Ɯ̗S%��+u�5Ʈ`�l��u.u�9���Ҧ�y��ڶ��֎q�8C�t���s3P��[v���U���6�ٺ���nka1SM3V��_��ִT	f΍��dڋU�H�-�sv��K���F�l�J�3�5q�FҸ�M��l��yP�䖆�Mw;^	�%I3�&��u��4��MŦ+vY���X�Z�)�f
f�a�뮒��.�e�.���j�4�l#�q��GI��L������M��	�Ԗh�l�p�)4k�jK��Vkq��L�A�؎t��
4Ψ`�R���Z�b\��K[y�g
	5�i���Wb���ˬ0f�;�4˓\]�-��-���m����l�<�[.VʹP������&�P�TMK�6̤���k�.
!,h�.6��ekKSS�Plm��V����n�H�D�[� !��ѫ��A��͢Z7Me]�ea�K3R�X�շmX�6g%ƴ�6�X���U�i �f�<ksNh]fζ�kA[d��q�؉�� E(\�0[v�[��.�v���e����sV Bh�@����k��M[.��6�s	M�!)1n�ٹ%�J����Yk����u�*hZ)T%--	����n��)1q�+�ڤ��.��]�30fd�%f@�5��Y�bs��na��.$p�In��9��B�惋v�����۔�YA-��B�f)�Ml�sqJJbjm1-�.M5Ivt�3f��F�٬�%�i3tAZ�f�����<B��c��7u?�x"���9���PIv7�
���G��(|�Z2��ҢU�Xz�p +�
@I$QM�T� J��B�	P$ P�!=��1��B
i+,��
H�AAa
I>�i$�&$,��a���}I (I��d�P�%H,�B�T��c&$2�T�(
DA@Pwq�BVI�`T
.o&"ɛ����,d1\CIěC4���6��l5��	�¤ݪ��6͢2f���&��svm
��xʘ�Z8�Qf2���y��,��eVa�����t˻���Z����&5!�37��d�**�+	QE�i����q5��Pr�)�2��E8��S��݋�f'v�����'��A�{���VQ;�I֭j��(/v��C-�l,�*.&0��L�i<�9����[d���)0�a�Y�a�RK�r r�;$���  jZK�bH���		��z=v��w��1�Lͥt�*f�VQ��ꗭ��GXnݏe �����1O,�1�i�֨ei��G���O5\�����K��;��N���'�^��y
=�rݹ�9���d�"1�Pxf���F��Vm�gi���t�Z͍�LO������BH��S��;C�O�;�e�����'i7k�ŷ~۾g�k}�|����}L򓹳g�.l֌b�`�
�f��gVd&�q2��љ�F��6嵔ڲ�]�cQ��6M����ؗk.Ьղ[���a��� ��!�F@%6��2��^a�.��a�LL�+.�%Ÿ�3�k��Fgi��mmE��m�ܩ��ki�S6+n��i��]�Z�ݫ����k�����4`PH��c��Z�*k-�k)�u�!$�q$��[���u-�k�Ͷ�]�r�,E;�d���sm%����i���ba�>��H��d)0:a��t�'{�4�竀�mۉ��f��*#�|6ki�Q�+�PW�=�뾺V,��;aU����Hq�� ��û�^;4�T��>�t��;�R�xy�9&2�zZ�=����J�a����j�e�C;|d��,��U��冽z�]9dsٲ�.�"G�O�t# #�P&���}6c�I��>�zG�V�eAe�Ñ�^�o��*��8������Z���vɶO9�s71:eKՙz�_1�}�m�������,<zq�ؚ`���N�o�޷EN������M�p�OL�hW�����Gձ�s����  kD�6����P)N��B�:�__��a�0"$暟��V �`�;�8#��&�J�>��z����H�3i������E$c���bP=m̖$	t�Jί�i7o���]�^Q�M($�#�b.jB}R�D F�"Ɉ�T8[5��Bܫ&}10�|�h��s�8���l�l���a������n���$8��pj�\G�	ľ�c��N�"ϝ�h�(��]<��$� �>@|1w�r`_���a{�"i��~4�����S� @� :��}on�H��n��z�N���^���J3Hv׿8�ٳ�7�o4��sZ|tm)�X-�΂&��Ɛț��a�^z���/T!���P����	�$�1-5;�y6������ݾz����tM��6ׯ��o\�_�&����Y0(_)0�[�m@p�U�}�8 ]OZ=���a`�7*�zaVne��	fQ?u�����ML1M���`B�č�w7�aJ����.�On����um��J�G.G2�ˑ5�.�d�#�m�ֺܘ��Ֆk�Mj�a��|��)'�[V� ��^ע~��L��4�QQ@CV�×~�.,�u��`��L�Ь��|��y�pn=����&	�ư��]]̝^�ā�s�8��/Kp��Կ	�L���'����b����t��Ȯ�L�`s�W1%D騬����&�F>l���}�ߪ��͊��G����c�AN3@(<*� U ��u��+�.W� %���>�Ǵl�x���I
��Xvm�\�{�桔SA��Რ��G��!�����\(a��u��j[0�32Pv�zU�a�X��v$�;�Ԙ��h��@���>�ъ��,Rst\ƨ���I���.M����c2|��K�k霪���V�vBp�B����v��T@@%�����Z)[ y|��>���������B2��_S	�.�A�q�D4�aq�6��P/%`���2L�l�m���9�����5q���\HS*��՘���3��W�auBǓ���Z�V��b��?�L��E0�m(3���j�|.������f>��7�/��i<��~�U��0�_�b[6+v�LX5j[/Yx �5�n棧�b_TF�� ���>&�W���0�=�����+�3k�/	�⍱K��;dfyh��&�#tK����[�����Sǖ^�^�����sQ�B'kɠI��+��+h��~? T�(K����	܊���d����f}A�$��M�{wᛃ`d�H�w7$d������C%�i�LB79qO��ʅe�����emt�H&�$F�h��!"�u�8�]\���"ة�rv6������k��W�v����Rr�Ԭ�G�Vn!���W>����)���P%�%e��T$5*ܬ��A]V�U�GV�]7��#��ߏ%�UNp��N�S������G�������P���s=�in�� E��ISZ�*�T�M��	��xg���Tf̧�f�^���1���Ĥg%�,��A7cc ���T�5ݼ�1���0h% ����1���U�ٽ0Um��&Դ�\��aVUk��mi�0�؂�>�c��}�Ѵ�:�=�/s��S৫�C}�g]��y֞����u�{|z=��"@-��	���I�^/��#(gH��Q?aaH�\�2~���H1#�> �ft�ʍV\�w<�C����t����o�$ 5A�����G�}��)���c=8�>'����m���y�o��9��9'��oV5����|�OI�`�@�BD ĭ����q�}!���d�N�?@����r�p}ev�E�(}��q��F��kL? �b�a�%'�$�|���vLM����;�Kƹ�0�eTx}րc�,}��`�F ����q�w���{f�'N=��=k�Ś?b"dF�]J�O#���]��O���<i�Į����S���8xBθ�@EM�$�?P���c=;��۽jb����@���{��G�D!B!ٍ$c;��2r����a["d��N$������cH��������`k�fQX�����x�]o�����q,>�^�F
RDP��L1!����1��E�b*�
 F�>��~�6\p�"}>�.�����u��^N��v E)�$E	 F2�sħ�1!�T mQ՛}��/���v�p�4�'�^��Q���"�������P�R�!@=}���u�t���� &'ӣo'�a�'D�ȓ��ߧI<����mEw{0���v��L{�8����(}"�H#��|��z�!��w���t:�_[�B����ׅ���n�HE�^�8�)��B�3b*�(�fLm@���/Ӑ���`��z$H�9;;n�z��Ϟ�|��&������6�=7�<�b@�þ�$��N����AɈ���M������""��F:���"|�7���>ӕ��!�p����iC�ƺI3ѐE_�#�O�p�f�Ek�LK?e�n#����p|~,�F�@4^nO��}�����f$�1^��gX�"�e
C7-�O���0���%�Ձs|��l�`���P9,7�e�L�%��u"}�P�m�=��"���J��ʨ����?�k�TY��Y$������Wj8���땓o����v�綆�H��K�Y-�/�ojkJ��՟Vbn_���}9���Z*�܃L����1��.���&՟'o�9��re�e=t"jȾ�;K\r15K< JQ^��_WVӢ�e�n��4��,�t�CA��V;6��T�q�6v�[4�-5K���6�Aհ�3IS+���=�7}<�	��"&����M��71�g��8�� =s5yˑ��.|7T꼵Q`��Tf�х�F;P��Q�A�c��ݥ:�z|�L��0�<�5�j����ފ"=�p�	�KS��F�.��i^gwVtp?w�;(��ks�A�mt�+$��`P�������.��M�;0	�#S��5F���+��Z�M��e�4J�
��pӢ�I�ɋj��+�^��E�ǹE�ŶAm,��f��T�-R��˻�~��x���u%�Jr-T�>��ʙ�CA�P��V���ǽ[H(������9�H����ƘQ#��!�7pի�3���2HJL5
3����`�$�w����y@8�p����:�4oŽTꂛ���r���"�ǻ���ΧQ��X�7�Xcc�ʻ=�8vHcanȅH��zy�i������I���}3qU�[�D4Z��R��f��TkP�A<����6�%P<�nI�t���[���P�f�N�{Q��v*�I��B ���4�bcR��[��v��ib�+t'_M��7�?8�SC[`F�l�����ܜ��6�qX�9n��*QX̢\���"��w7�GJ0�3! K�)e�#!����řG���ŪN���e�8V�+꘽+Q��`���7 �Z�Q�XL]��G�i-��*��h)�s6�@�7E���ų[*�7M��������p\�5ցb,[����K4�젢���ˊ�_���sCA�\��Pj�Rk��%��1���:mr�m]���:;n���6@6�%u
[v�F5��A��h����m���RWr멵Y��M�����Y���1���l�v1l�ժR�3�Ѳ۩]R�J�����d��R�ypjg���2@ k��mZ4��.�]n�"4���ζeIQ��%�`Q�%՚�e�[�XF���M���-1�I���3^�*g��q{0�F9D��6����*����"'(���.:�tg��ι����9�Ao��nf�Q&3˺Q4����.g�"0!��I8��+G�N�x^�t�#f���Bcz���u-���G��S�u1�=-oq/����d������kҾ��H�w&���j.}i]�i��}�2��� ������#���n�I�ǱB\`>��~����_i�8�z�FWu�X�r�1��Y���{�J��uB�޼r΍ހ%���W�����"���n��rM��J�8*|�f�f(�J���ԯ ����qTrƺ�����4u�������S�9!�w{_5wj�����칌�f����+� �p���J��4%BT��U�0u�/�!�P����/	��S�rI(U7��wH�*�*qޗ�S����!���nu(�9��m��1p��T6mԒ�@�׍�e:c��F񂇡�����μ����}\�� [�P�Kcc5�ن�.N<R:K�����G�Ye�0���l�\&��K¸�����=�g ����PxPV�ɍ�A���uU��8g�唗��2rޜy�cܯ!뭓���&�V�^�]���Ӄ� ;�pXm4/�S,�>�W�N[[f{;��>40Txͧn�y��b��_t��7��ȺF�e�����kcv��vE�U�ڰB�o#	J�t��ǔn���>H��z��D������C��̨E��7Y
t��0��L��w�xz*��^4	����D.��{���0��n'�OO�0�h��/�TDO�ߙ���T=0	����{�yS�M���1��:�1P��A�!����룛s�jr��T��w��s�j�#�Tz=Sw}�a��2�@�E�2�Wՙ�l�cګ[i��q����'�m�c�;޹��9�J2l��x�\-��#	����Ǒ�����ox�ne�D�@ű�:ڙ
Ol�-�J��}���,3�$<���p�����w
z��b�r��y�<`*d���E�[�7Z�s��
㯇���RT��qO�E�y)���rݫ�-�Xfb9Y��0,-5�m�k,��T��DV�t��+f�����s:2UYٝ��^�vzUT�` [z:y�s�i�	�y�LY�����e�ӂ�]��u�2��9����]YFQ�@8,��(%�P�r�3T£2߆uT�ZF$�ÌM�(��aG���\�|�ɼ�&�E_Fb�p>�=�Nk�30���h��[dë�r�����~�랎��s�e���h&�>�����:X�:V=Uw�gƦ��J6�r~�pZ��Jc0򲾉�7�ہ�ࢲ��"%͘UK�%��1�Q2gaD�����E�CקaF����hf�r�yZ��8Nm�*��2��qc.�H�^�6�����)�saBmL={QD�2��R_n ��&�lҹ[A�qn�M����b�H�� <����|}�Wz9B[��i�^Ѥ�p�ۍ��~��H�9�6�xp�I{�ќ`��a	�a����I�(P�Vc�%z�*��3��9����R�^�Uf¬Fa�:7��0&��j�N��ӳ�R`�BB�ú�Y'�r�l�}h{�9����D�v��eBY	|�aCjoB@�����EE[u��[����?m��e �)ʵ�F�]O���y�nT{�ѱ�o��`�Yԡ�z��]ї�%/1�=�PtM���oƐ;�ߪ2���J�R�-L��kM��:0�t�]�r��8��C<J��Ç1�f�U_�5wMF���C��7N�f��w��������c����v�{�cnߡ�7��7Ԧa3E�h��F߯���W��(A����3�[�ݪ����bn iǻ�<�7�(v��#��=���^��oU���&��t_��>�X��k����{�3�(��OT�@Fk;B�}h�����ҳ*2H[XQ@{Ǖ_Fe�~ˍ���շ�|*E�I�:�I|&����O0�y�'�)^8�B ��b<g��P���l8�
x��ۙ�ѱ��LG��J�=��S}>��g;��z݅�$6]Mj�����EB��b��I��,2f@��᚝�S+i.}�vE(�$�ug^\Q��V�M�{�}��@]t�n'����*S�/�D��S$�rb����þ�C�n*fKYY��b�� j;��7Cdi�W�ɻ�����=��u�}�%�]	K�Q>������w�53[�/sqM�_+����n�s�k3Т]�P�37�ݗ�5Wu���Z�q@)�G贠5�̱���#�dn��)cc�]�f��l��"�g�L�[E��6�Ĩ(���'����ֿb���&�'ub=>��sM�P|�{D�}R�`WҨ`U>�d��:�H�ף�"�.gH��)�G��pZE����{/>lu{\��h�ʹ&=���_���L���9��s�5Ho#$���-i5���'�}��q��05�Ny�T4T3�~�z}��P�	 �j��l0��ٜ��s3.�_YB�.�_Gt�w~ܩ��]�ۓS1���X�S&�1�a��Wֳ!�����׵vdI5�L</�7a_��G����.(J�[%2�r���$�����M��A{�f&O��:������ʽ�z�fe�]��E�J��1c�n��5;<�s O���N{�TH��T��<�am�JN M2�cu�uW��R�pUVI
|>��^� �Ƚs׎�� ^�L~Hj9^Ǝ,��U����ԭs��=�+O){
�W����$t���O���d_噏�;�|~~���I�6揙ϑ����3�Y�k|�<�ɭ�,mmTV��LfH�L=�����f���;ڷH\2f�\MeVF��skջ�ҽx*�K�zS�بW5��4b��R�`e���W[�hX�{�a�]����Jn��K7N-o	��N��[z陕�f.���ڤ����MTõ�LV]��2����]fl��͘Q�&CgR�"A��p^��4�f4%�e�(���S��[)�tM�X;X�Yl�آ�[���Me�5а��.M]D�g6�S���ť!x�Zl%v7+.u%���9t��\Z�K��m�L�R��.5�8�K�v4��8�f�� f���NprBu�|��mI��[���s.�0֐�[�)�D]*[Kl4K���a�m�T�Th����\�$�5��77��wO���lX�o�J���j���bS��8�j�\�;�Y�k��O��6�*��q<�W5����[R�E�ه�J�s;�9�0!�H���+zU]S7A�S�F*����WF��,D�b
���垟��L��k+e8�]ў�V�U���w�K�a�~��*h{v��ߓ��Qn����S�PYE�`�i��᡿E�۽�i"K�5�Pq�r���8�=���T�p~\�9���
ϥXcl{��O1�������ۢ�:�ɠ/۬���L� �����P�l2�b.ocA4y��{��"#��|��=�$]�Y�G����0j^���^]ًڲ�5ל!�d�ST۫"����~�]�9(,b��^t�N7�0'��-�R)5��Ў�M%����<�{|<'�Ew�r�;5E���t�7��Gt�2|�f���Ϫvd�2��s���SJ�������ˇu)����@?@ϒ�	l3L�;Z݂S[.����3�rƬuJ����]�L&NL6lmh�>Y�D����w4&
���o��n/
'��$�V�	�F�5�(�"�)tWk���x�vf���^�aT�S4�Ow�.
@���!��l���˗{���_,�Dx��3 @`4��������tp�P�*TI�3�P�xnF�U�|˸��t�+���S����Mq�^U�J���Qp�M�w�OM]�eTM�D�z�%�`�7ޮC�w��8�ד�@Pz�gn��ϟUI�]�n��S��WY7U�tn���S��۩��o2�!��)��I�tWzs&�\���z�3��Ʋ�[fx��R����y��qy�[�T��Wa����jl�~��n�����w�����r.������\?��ڬ�3ꚨ���>-fwm�pG<W��#��W:�q�V��PN��y^��v���g>쟹����6��TIY���Y����7\W)�[U�x�E�~P@�p�&I A�6ФDn҆�mA��҅��շ$ل+�S�����]���֝ec̜���x�>���Ǩ�J�bb\ʬw��Tl5��P��n�v.�w}"�$��*�S���n�õ2q�r7 ��i�.���Ωeum�M�4�/�:2����ċ�A�r/���NgfpO�Ѿ9ʷ��7��9^�� Xb��v��[ӗ�wI��MheL�\}�҆�M�(cx	׾6l���%qk�lc��0�ưx�A��
��d�[*Y�]�������_���!��@?ګ��a3�~������~����Ȁ���H��n���Aia+vV#��d�*vr�Q5��S;�0��p�f���L��7cfT��G�$\�\��Lцaˉ7�ifDlj���(��B*�(sqe�ൄ����mFk��)��0фn�Qa��Pk��B>��*��������>�[|�r����,�Z����^q+�	向MI6�$j��T����;�~�a{�y�\m���AD[mg��ԩ\L0+��ܢxw���&���M��*s��+��mQ�m�����g�����j=��1-�>�<0Ã	�AQ�r�3�q/j�_���%)���P�u�8�5�_�dn[��{����=�)���x���[��i��*�ٞ'�+cw��5.@��z��ν|����lke�k]B�iq1]+-Ѯ�(F룛a�^B7gB�ˣ3\��w�T�xB�\��j�m�Q�d�+�C�^�ژ�7O|k���U�vsR��ۿ{f3����=y/5/H3��R
h�� ���Ʋ{u���ƥ`r�:�t|�5e��K�'y�ʫ�<Po�:�tU����mjR2+-�r}�y���:!y۴t�}^�rn3�I �%�X�{���~�*�[�W9�U2\����3�<�Ѯ����J��c�����Ϡ�ڹ�m0zseH��4#�8{EW�C8���
&���pȅ�T]q�3���-�ﶭ�?]eU�o0�|�Ud�= �l3�vA:��6�=�����᠕i�P�(B�|&*����=�^תB���*�=
���Q� ��"غXn��Ec{ڕ���iBp��ߑ����1K;R��N�Ä�uyY�䤋���̯u�qj�%ꗶ_�����������d�H!m>?YH��"P,Í]�j��h:�Li�pn0-�ѷd�ܴ,ͶV��Ī�������<L/M�t��r���uH�*���o7e����y��=ǌr����ueA��u��R]+�Y̼��y�4O��2���r����G<V��W�siz(������ �;�e-1��B��̜���P�A�':�$Y���^�V=F<s���D�D������k{F|Y�6ϱ�X�k�T����w��N}m�71�^����^��<��5|b\\��=��+S�tf�Oyt���`�i6�g�1����JC}�ڼ�͢���ݫ�r_�u���0�<+afFx?.�gn1������U	�8�+�.'�P��̘�3��Va6M�Km���m�S��׮����8�`�2�i��/ۆ��D�+���������7'�W�׸��d^�W�E�X�g{w?_�������u��s����=����V��c���y�����ąF����i4��]E@s52MYba?��+(ʪ1QWk��� T�,]]6`��U���)m�$`;B��h�h�q�s�0^2��*�P�ܵ�Q�ز�E���B��"ڜ�+n�Zs�v`���"�"Z[P��>�u�8�n��%
�	��.-��0ۀ[���e�-[����[vLMPq3iH�Ce�v�VY��v�U�2�f��+5k��aK�� ؔ#b��ԅ0��ml�Hr�d��h@6%���[)s�K,��E��[͖gsf�r����F�Ll�t�m�L!ACh�;&�i.�H���k�U��n��gq�G��v&�,9��.]��r�+:��t�M6���aWAP]�G:5ΔZ���ꦤ[�*4�%�Ԃʦ�p��W�{�f�e^F$�o8-��-~�{��7gj�\�n�/	��x�%�3M�2r��N���V�&��[���L��)j�a��`����h��ܱ�P]�Gsc�<1:�	ɨ7���%X�ig��/�9L�d+wt����I���`��=�r�W�k�O a�I�<�q�̈l���T��X;��/ܞ��xAwn�~���f̬u�������j^�wYH&D�2`H����jY�����K�������@�R��>ۧ+T�Z��85�e&Ie�B��Y-�'C ������ۊ����Ž;�ޮx+}�vK�h�uM(G�Ꮎ��@�eg��TW�ÿ%����P{FM�E�RB. p�����>븧7C���j�Rr���Ռ�8w���z��%X3*g���7��CC�Pw�O��w�M�6}22�;k Q��f�c�hL�"]�MƷK�h��^f±�6�ǚ��[�]�˶��j�h�,�� C�����q�Vñޤ�/�˧c=g��hN�q�	�y�7;݈-�|∸��j�}������r�pG���:�(��I6��w�^ku��������S�W�>Q��G{(��0�rQ�q��T=y��Ȼe_"_1cѸ}�k^f�R��5�Ę�.�Y�.���w\2�v,���hxE��9Z��Jj=�����~~Rڧ�&l{�����wWwkK�d)wa��ȹ鼋��8��#�E�R�ڄҌa��N��-���G0�zz;\]np)�W�\��w>ډ��l�
������V��u�@��L/����x�����ɘҵք;���@�@�`�=5��u�f=kqqΊI�X'Щ��Sշ�� �')�g��>8�x�>�~v���çF���6
݊�>����YV+Nd��w�A�3�����Ք�B-���<*S9�4ů5[o&�3�]���kmԳB�6j1A��u�Z]/�)��x�j��u�����S0�R��٩G����[��Ӟ�[׋.���O��f��
ּ�Ϻl�A����)���!6�}GwԈN�v��ߺ*���<��̈́%C��H��>�t��q�M��K���0�y��� �	��G�*����	T�Nyt�4e��umS|���2��wC�~hD�1t/���4o�N_��߼�q����3uC�ړ2�8v�LՉ�֭Ѩ�ǤUU�-�%+��m/M������!��]���%����F٩�;�-��1X]�T^�"�=7U��l�hٱ�*0�	��.��H��`��3�¦�z�G�2lљވ�ײ�Fg�Oo'0:��S��{xv�ɧ���Ꙇ*AG�B-(m�`��p�N��*xzԋ��v�M2�dV.�r�%�==V0��^����������7�ׅXa���9N�֥��sE8J{=��}��������t�����,��r�8D�v��)�/Mc8��C�=yJ���p��]S�95^��^�|OL�mI��m^I�ߙ�e��d���͚EH%�ң��&�9���P�0��%�A	�2�d3�(H�Iǳ�k���]�K3�I jj��W�i�we­0�]���#�F���K�WY�y�Ï>0�s6���y�	��L�	�(�����y�x���8 ���Ç�~ZW��Y{��vy1���3�yvG�9,���y˼���8G{T�*XvUU�z)�^��pXd��2�FM���
��<,���U����ٙ��ίRWr}�<�b�DSoՏ�ۜg�ao���$N������j�1�9L�$�>�_q'��b4pq�����-�b��V���h�BG��c1�1�c��w^9fz�-'��/��wOc���]V�U���\#p��E?S�k-df�)M��l"[%8l6���[��/��uͷ>�d��}8(��Ċ�׆�'�U�����5��{=|�Q��KT��N��9�٫�n��d*Ӣ��B��D��E��.�����[�An���<ыDv�-٣H�5����5�k܏#��+�M
3>�q���ƗwT>U#ѷ��y|��HE9N���=�9,�՞pz=�z�_��z(]H/��`L�u��rh*���g	c�5EU`�� �U�Ol�s�ƪ�=~[��jϓA@9�'/��R��^e+��0F�-)�w���(�p�iH��>A�����z�6��]~�8�M7^/k�zP���㐥�@gՆ`X���P���-^4�t����9h�t2������vge�1FK��m �5���S�mK�&P�^H��r���/��t������0�/9��[��Y^��������ŵ;�����k5��V;���¸Ci4!0Rqd\�L��.�jע�_L�55\�êȬ���/�e�`����v����!�Xۨyqjֶ!=�qs�A��EY�E�UV�$N����$}���/f��b�����{�X*6�7ȁJ�F�f�	�]���.�a`���\͘ۉ�EK;n^`��3n�$¶�4����sZ��5g�ps-�[5,��x�Z���Kjb�ɽ՗l-9sFT*[�a�Y����ғ������Yr�WZZKr9V��l2F\�4�]�R�F�u5Ͱѷd��b�l#+�6�L�@Պ�b�xA� X�i����x\��lJE	�*62]UF�7[\�Ŕp�ɥ؄շMR�]]Xf�vΡx�]����MtuQ����Y�t4(mV.-�]���i�TWl Vh!,�V�&��Z�����1D�������<Y�,��-�mˆ16�<6e��:j\cX 7�#��l�Z��	"B�p\&�p�����u/�6%����{�FzFv�Z���|�cβ��-]d��K�]�����z�ܭ��WQ�b;j&�=��mEd�d��G��`H
`���"���ÖS�&�ۛY7+\��S^�_)wV.�a4��7�T��>�T=O
��g�;wW|�'=Yg��oyb�Ѧ�q{�=�"p�M���8�	���w��D������{V߂��U�b��7���ǽd�^�'��<tf���N3D*����9f�MW�d��7���0Zf�O��O���~6����c�(�	{���ٸ���s��K3=}4�69`!Gr\d{	 �h=*����5�7���I8>338�T�k%W�x�P�^uMIL��q�*�K����Y�����]ls��V��'l{�o�?LǭrV����"F�L�Kn�΄��ˣ�9�j䍵!�0�l��+4rvN�r��Pa�~���fJ�L^��_z���q�R���U�w���K�|�W;�Բ`up����V���k��]1����l�m⳧+�Yr{gopW\^�=мŪ2��DLIjI�������S�B�m�D�9#eD�Nݞ���6_DאM�Ys1&�VT2���8-���6olL�O�������4�=yݽ��띌=��ۊŃ��5D���X�9�.S,��W�����$��Ysp�P���0�d@m� I���g��}IzjL��ts�-��;=�)�^c&�\'���q�E�%��ʦr���S���:³�������QM��;�
�N$z|����W�����Z�@�y�Oj���g��Ty�q��1Lgd:n�ʋv}��^
�����O�kW�s�����"DB�f����ci��p۬K���6�+�mu�[��¢��Av�0[H8-��eÄ�m�ov^��:WeȎ�q+������T���Ə���j�g��1(�Wnz�߮��<�o�����O3PƠ�&� Z9�ר,���ޭ��ߛ�υ�rWN�t;y������(c�Y�ں�[�8����A�7|��}q��fgN�i�BjL0� (h�KO��yNyD�+�:�W��f{�[�{��ދ�Ȼ�'��4�Lʅ7VDc��&D,�>�tl�r�#"�{ ��/4�3��4��8�sB�V6h3$(����9�h�(����Wו�!�'��U�2(���cV
d�e��̸�^P�����w?���j��E}�#��;�d���Ꮥ�m���n�-y��۱�y�-Li���G�i6��b��֧É�m�y�VZ���VJ���k=q���wn�q:�w-�C(*���S�dg��"NӍKdzpVߺ�:�.�/�!*�v�B6ZO�W���w�aw�>[M��� �����yǦ.��>U�1��1�O!���ɩb�O�՝Ύ�[�q�f;D� 7��oH+m�٫���&r5�ܹ���Z:[���d���	l���m�l���߫�z��;���q�vUz\mQr��3#g�I�w�G2bqx)�k�'cTmn�x�wj�>�'T��`C!�p�NN3���x�ET��1B5gv�L�4��#ls��:�(��=[:����&*`��\�.�j'(y^FU�.R��f�{��jj
m"�B.�^��Y����Q�+U�F��x(�O����B�s�����8vFx�L�9/u_b���5{���y��q�fS�Q��#l�Ӏ�E4w65ޕ�r�)�h����m����yx�[+�/��i�}����
�>�i���fh't�	�{�*��^�����4x�� 4Z%2^)���g�HKLP�~;���+�����ǖyܜo��!G�[U�ꪙ)7�Qs{�w]�k��B�^��F�P�Y�F��S������8��c4Ʋ�H���0�W[f���&ڷee�
@7�N��3y~��Ss:j��w�%F����9u�ηkZ�����3���+
�q/�`�Zf=5�/%����+e&-�Y)���`^^�T��`캎���s�U����Լ�v�0���������7�{5��`�ݓ�a�I\�h��	���M����
�鮊5C��T�neia�u���B�� z�C-\��Qp�ч(#b��n0�W�������r'V������jY�gF
���L$�i��I���۝�^�J�i��ݔ�_gtI*�������!��;��c��T=�o<[[�d�'];�^Z6&%9�ē���n�u����X�� B`��h�	��5��`��ܠ��n�OY�R�V�`�sH���4��3���<��yngf�W��7��/���� @D_�UI HR�x�������Z�`oy����qqa�B�I#����}��!	;�BI m��H *�����Bm���Hӻd	2�@?���k�@�� ��Bi�@!4�			0����ў_����a���n�M�� �(H
�7@�4�5�)���C����΁��A}?L�tC��Lv	�q3�#�	w��
�lx��.UL��ݾ^A�����?2F3�E1XH0��gk��0J���p[�˟��n2(w�V�K�T�A�����X��S��	�}�m���$"������IG�⸙������N"��UѾ�b6�k7���	�!�i���J{gZ���~ñ|!�{(ss�����=V�A�c�ÒU�V�$&���]J�F@ش�}ګ�q��q�;�`KOl⁐)�sY�_�o��[ ��P�K1Y��z�;��>?s�_�О�	�BKkD�PUE`@� D���DTiDD��4�AT�b�E����(�`2�BL���i�t=uC�^+(Y�B����F��҅��h��sc���P�������=08J0���>/C���C�!7i���
1��(
;�
�������fI�w|�7r���,��+��E�*�n�,p�K������A&u�|��׏�.�6�*
j�3n��,�?�!�����u�22�bh�E����� �U�QPS��/܆�&��^�Î���T5BXp����RHInn_uDa��	~�Q9<H@��'�8�ɳ�w�2C�8	�Gԥib�agٸOi<Λ��f�\C�3�����@R�hD��p�����˓j����E��tkBY�]F����{����K��GA���S�ǔ�?ô��N���q�E��EAIǣ�C�!YD:M�8l	E(���\|;���}{����5�� ��5���8J4.ai�5���F4q������ٟJ~Xv3���I����Z9���B��K/5��\h�7\����	�dVKXns/8
'h�i(�^����h�К��h&��
�#;�%*8s��q�f��Q?��tt���3*#��Ձy���1���)P���������7��C�md;
P�1]>�WXh��ܑN$)���