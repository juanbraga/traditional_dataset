BZh91AY&SY��e �߀Py����߰����`�|>�x/�Cϫ�
:�$��0����Ɉj���10h�S�R=&S&�`L`LC  ���T=@4� �  hh�  S�'��OE�#@ ���4 H����4   @4dhDB
zhMO�ʞj���6������4&����HT�*�Gp@��X�t?n�~@!C*A(p��?5
�Xch��G-�{��:���˭.����3��ȇ�2A1��l�}�$�$�o��Z�]�;��p�|�h�(Ӥ)dcIM�5�L��#+N��'%�,Ē�"@L�3��pm�΀̥`��ac���9�c���A�Gl(Al.��K�ڶ�\3��q
C�n_�YXC02f���8^��l�hޒ�$9uP�F��Da����- �M��dZ�B�j���ʡ+h��:�i�,&2/p)�q��#id���.�꠻�N�hZ$>���	#|�U��m�Y)��tƪ�_w�$�e'��jE�iDûa�!��vE:J:�L��5��+hu"'�ظN��=0
�����{B�obk�%����
 H��
-@���HRAPcVd0�d �R��0���wsU��-O0K���s8rG(n�����cU'��,�-ɜ�jk-����H�r�L�Z���(|.Z�'�"��&�
	�W�Bԋ�h��x*�B��K���Ihr�4[-��k%؞��R���e|Ihō�B$%�whÛ�ݔ͎+G��[J��?O\�I�H�hIS���	��(M��d���5K�b��!
���|�`���	�!gD`���`�m@�I��4C�\b�j��gĀf��c������/�5�@v\���({d����
�r��,��Ɇ��e��3�6��U�Y����D4�8�6]v�\\A��eD�>����Yw\����'a�ԋ`��S(!d�o�A�[*\�[�Z,�BSl[�T/+�^#	n�tsH�_�X��yI[���Sj��T0�X>�Ǣg���0��o�)���V�z��=����r��1�HL �h�I>�:����}'r1V)� �Hqz�n~R<R���F����z��Uy=��w��ʄ[�}V��<D��s=kNO�(��oņ-��v����A�mڏ���t�-CzBp�3��5�n���������*DxMk��^B2:�@��I����X�9�	�am=�@(�X�WXU=$⬪U#�p����(���S�Ͼ.5A�j������
J��D�c֪�H�PN�����Cc\e��$q�]F¡R49㤟~0�斀��K��py�7��%��g��fLWc�R6n����>3j� D.�Zlcw��n�3E�hUcX�"<�v����A��n�<�g~�[���!�2�C�m[8���$Pգ"^�M)ij&f\��/� �n�1�!�W92,��@�+���9F�T��S��L+q�e�-P��ɌY�ɐi�Ω���H�
��