BZh91AY&SYͯG� �_�Px����߰����P8I��Q �A	"i�z�*~�����Dz��=OS�hѠ��Sѡ��@�   4 �ȈF���47�h�   ��b�LFCC �#��@���oT��4�!�F�0�z�][Q\AK )H!� P���?/Eߌ2����ji캀j �P�>�^�e#մ�����tl�B�R��D�ӑ�Kr��H��q8h�6-]O����w�oE&�h3d�XS��e�7��`��&�����O�>q�r�Dg}��I�92D-b5�ec9{;�g�cA ���g�Wt����_�:�?���Њ��N[o<����̿�xf�+nh�s�Gۋ�lw��_.��4��K�$2��yF��j]�][]��)�	CY&r�4�=XPVASX y��������Ln�|Ϋ@���\K��qu��Y�/:�"q)K����e�b��=�����g�['i���D���6�����vM	�Zε2#{�W�v$CLn>�%
Na�2�vc���87��|�8��5���ٞ�oZ3�����أ��,�:c͜�Rkg�n4�nV�ҁ���OVȫ���S!���T����$�Bb'�!:�/7lFAn���ިd��@�w!�[J��'�%��Q�	�6���B��ؽ:��*e.��0��k�O���Z��3�����Zo���_�&F~�~1 �7���8�}:/?~a앝�k>m�ySf���9/T���猤Dj���Wmg�.��Y��z	����l����z|i�b$��eH���c�w�>ǹƗ^B�EW��E�4�k_��Y���6����I
�y�?~�{�1d�� �)Aw�`A2 �}E'O���1�������D-Tә�~�p���t6Q8�-�$��6��",�f��icU�?���L��GQ��0h�&Q�R[[�w���K�z�$�d����s
�΢<��|\�[2L�)H�@&9֝J�o�2����)��K�J�iP�Z����ey#as��"Bբ��%y�HV�̘l)hn?�t���Bb�&6k/uy�ؒwj�+�1��{7;B�œ#��/)t���rID�qf�� �����B�}���$l�4��k^r��f�P[&��4�L�ZL�᧝B^���$���&�.I.���a�����I�GĂVۯOݴfՓ �:8��8:^Q�u�GyJN��mzC��P���<���Q�tk/J��PYz��&ۆD��D"��[JYY�E��N�"��L����T-���]���Xjwq�D��2p�nZP��_]5�g��5�!V�
���4"�W-��Knu��V+��k�׌nfG�ԥC������C��Y	�{�Šj��"�(Hfף� 