BZh91AY&SY��E> _�Px����߰����P^s�`#��ca�O	$�#&�z2�jf�#iFM�4*h@���  � %=D��SL��l�3H�h    s F	�0M`�L$I���l��zi=Fi4�=CF�h�G��@B�P��hE$�
�J�Yп�g�HڀL�[N�pu����l	f���/.}>��`L���,��I��-T���J}�p_��p�.r4�D�:��j��.��%��6�o0��B�1�����pI��m�k���`V��+�x�!+lƉ$��xw�4_��8��f#fӧ��M�7~�C��-�vh�U9�#�;pix<�`T��c�p�o��t�����@| �RX���eh��
�-�`LKd�� �a2����N�86쯘����D��0uҝe�Z�a�3�6[+ �זF'/,��UuN[_T���Z*�(��*',bs���kzGb�aX�����@DSX�ʋ䛆���P�[�cE6���S�jE[#à���|oW�PHdJ���V�#�Yb�a5�mWK;nUH^�F8�(�X&	$��1�`�0�Uʛ�7 �%���%eR�$
��c$���-6�yh�u�����p�����ݐ���>��u�F�]x�wx�U�.ǷW��i�i�ߵ��J�ǪC��q�5m�S�x���SȦ�m �!�B�s9���qD�M��(��x��ҼF0�Ҁ[��7#Ｄ����H�!sܕ�������EҢ�۞�tc�p�f/[jY��۴�u� ��UB��^�z�e��-t��@�]��?p�BM�3�UѾ�P�s ε�\C6��a�"B"bE�r|�R�M�+4
GsN�T���6������ i*vtᨪ��C:L��;ص����]�����Mٍ�eIC� ��Oa	k-94)�%i:��+4��	D�H��8/�%E�%(-�e�ΈP�,K�$����D�J���F�<��!*k��f�sEKw�P�Z9� �^�*)�?��7�>Q��_��6����#�{;e� ���
G�85����5�9I@��]�2"�\�)XeJE��$z{Vu`_%��N��^N���IF�����Bw�,�*��q�Z�xޕd��5{3�XW4��<hy&[("�F��Y�J����N�5�\�W9-qס T̹L�vg���ld�j��J�NB�H�
ȧ�