BZh91AY&SY�ڠ �߀Px����������`�}Ͼ�Wf� +�3f*#l	$M44
l(Ȟ�i����@� =!��P �F@i�� T�L��    @ OJH�@�    �"�z���� 4   ɠ	�MOj��<��Bi=C�M 4��!��"!j�@�
�2�%�$X�v�j'�uMX�LHC0��fC(I#U����
�v�5����[�P
 �<�p�2C����ݓWuܺ��Rnq�8����?��΋�JR`���'a��^�B�<�,�&T>2h����(�DQ`�$5&HHPM[ �x�7i[�RU����2�
��A�dR)�����tё2�q�hJe�y���m5��Hez���¾Hf��:s1��T���W���I��HjG� 뭳�<iL�H�{g��w�E�2�av�y��U�YUY5�wkakaIO0¸W	�x�[�@�h�.)�9�����ѓ�bYB�#,J������e�w,�mv\v���M2��6Ǩ�c$� �|a�K��x��Kc�4�������R�\�U:/4EZWo�زU��&Lv#d�;�l���Y�����61�+�Z�`�o����7�w{��ug���Z� I��&�\�"���Ƀ:L0,��i�,֡;�;6C阡ŷo	.!�ё�vۥ]t���f].�.�֮P�,H��X!��pv��ė2$!P�&y�_Y�24���E�<k���9��0V��s�w�};��@ 
$�;S:i���U95׌�"����:��l�b2Rv�)�U;RM��� {�C��0fh[�/�[x�7�>�x�5��2��,v{Ln���L"v᲋��n�!t�o8��AS���+�x&b��Ba��ޛAe��55�h�]¤����+�}���6��)�r]趇i,�w_�&��	=���%��� aWHTu�4�x��^"��:�ӊ�:���&	&��A����GL҄�y#h��ӫ5��C�N��l�BB�ʜ�����کX�a��Z@ |�m� p3�?���)�h`s�⨧b�S�H�$�E�J��%v
�$�0i�DV�AD� )'"$	�m6��B!	���J$BD��$CT�\�
$&(,5��3g&B�"�C(h^،� �b�:���4z
'��2෬���{���;����ї÷�9aWe��r�O	�vY��M2�/���w���v��}��1�c�?m�5�w��R� ��C�L+��w�ja�^�Q��>f!e��5�Q{=�������ې�p�6��cVi-6 O������l�Y�\�ԇ�C4��6�=0����k����S2t�=��iF&}�%e�(d!滋�����lP�D4�bJ�Q�5	җ����ULQ����P�M$h �U�暸f[�>
�B�@��J��TX��%��HED<˓�ӇȘr8�@��8�InP�tq��۷�� ;���=)�ʲ�c�R`g2����b��]���`�D�L3&����כ�>n��<�k6H���'�I mh^E��r1ci͔0�b�$T�%	t�E�K[lcDQ$�L��BA �T�yk$qD���' �\" �,
+8���%0��TI�;ʊ�+P@c�fm�BF��%��������ۨ���Ɔ��W�8o��M��A���JE�sy�z���ж��Ga�ݛ�ƀ@�e��2N��7.A��H��x��с�T�3Ki�v�խY�PO��
Q�M�}���ه�e���D�V�}��Rne.�uO]���9�U�!ⴆ=&j5#SP��B�<��.�)I��}7�L����w��������V�}JKS���]�E���1P�wc�َWJ��u�n^m���H�
�T�