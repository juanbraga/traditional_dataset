BZh91AY&SY� �� ��_�px����߰����``���t AJ�R�|       [a�+G@  �
��ي�� �h�E$# ��d����"�-&mP��ٮ 
�%�� �R��͕T�����`j�Q1����jH�iJ���� 6��*�f�JJJ�i*J��J��R�DS���)Pd�&M0��C�*~i�����       �L�1�2`� 4a��H�R�� �0 	�0)L&����?T�*<5O�=&�C�4h3Q�I��&JzcH�OD�F��i�H���:s��M4��(?=h�(g�$ IA�	@���~��q?4�
,	��@$)�}����`�@�C�$)��L2�	!L8g����G��c��@� ,$XM��AdP��B�HR@=) Id�y2@)����2����a��
H�I$"�,"�E��!$�J@H���)�H�B���r��(�����3>G���Kv�(�|]f�����P*�6���ɷ����0�Tf�0g�j�<;F�ЬV=��d�{*[s��@Uw*"K�Y�W��cS5�-�6Sn�Y�&�Lպ.@�20�ȕ�2�e�BT�՜�iM������H��T�n�J̃v�V%�.�(���L��SJ@ �eڬ9�ދ�o.�l�1.-E3%�c�Fe&�J�L]�F���i�R�XU�R̺%����f4�)aX��2,ݲ��{���e=�?'�2:e�NLw������e�yx(]1V�{�R�%8j� �H���J���+Ā�m�%�3ݽ�����L�a
w��t�qDdY�����*%���f��4�4��$EG	K\U�%�Y7M"�U�X��r�̧����+/@���n�텸�ˑ]���i�B���T���ژ#l�$�V-n�F�&�	E��Ǉ$?���0�b�x�7R�]�����z �q�����fT�,�]%W�GktQ���[m�Ff��xS�p]G�%��7y{C��b��H�X.n�u�H�ʋN`�Sl���j�M`���c�HVU�@�Ƌ{@�+m��c1�m���[l5�&��dFB��D`!	�.,!WmnIggt�l�xh3
ӄe�r��"�&l�;oK���:��AZ����4��mn)���#弥&;���-�́*�N�+ݡf��\۫���؁?���F��],�䯆!��dP�Y?Q%eHi�p[0�[f��F�F��F�5t����N��͸�E��I�fӏ����re�g&�m�a5��$�Z�I0��x`�pk�w"���!�D��[��E��P��0ŗLF'Jˬ�
�$Y�(c�A�2��zX��[twNi�x�N؄���
��cx����-5E6Yy�h��
ú�Ŧ�q�׀���載�=�-�i?�s$��j1�mTĖ���I��!8c&��9H2�!�/M��rfS���V���U���7E�L�v�3&en�[��-�KۢŦ��>MܨuF�ub\�p��4ƕYt�k+q��t�^(� Z�YxjG�.�f����^
�n���&�Rn�VN+eM�(� �	M05�
b�����?���+&;���#_�Q����x߅�&�5�&�\�t�)�0�11]YD��Ck�k��5f�hĎXClÍ+u�� Lm5C`�҄q-�i�0�p$k�E�Y���s�� u�Le�$&Kr�e)12JJh�J�E��L����M���6�+��rF��m�CE��)-�l2�-/4s0]�z�v(B)D�SZm	h�In0C�|o��=n[x,`S���nH��]�Y�U6��2���j�1Mm��an��2���a5ֲ����[\]Ki�\^�QK���<�]5��"Ys͚:����
S.`��qJ��ݴ3�s��%�+h����u�.�ҖQ�h��4��˛���̙v���L	1�씙
X���6ikR.'#m�0ۗKQ� ��c(m)L����Q#�WJ:�͖�6x���ƉԄZ:�P�g#�eY���ĳԖ6�b�]eB�I�%k�J�nC^u��q)�k���`t�`��%������`[ ��]]2�L�D���e�8�k�[%�H���ʻmB4�;L�bU����5��1e�Z�a��qe�Zl�)uځl״�ͭ��A��3MT��H�U�3+-��Mm�[ͻ��i|�h����m��]j�4��ڲ�JM��])��-66�F�pF]�3jj���I�`�f56�-6R	��e��3].���n�%�e��nյ�������LF��LJ��hu�f;L6mi5��,��ۚKcĺY��L+h[�ݢ�]�e�e/g���pWe�cZ�cq6�53�F�6�v+lV��)�3.�-r��]�n�66ٕ:�tV.���1�7������I	p�t��d B@�}��B�����B) @$X@FI$�O��>�	 �Q�^S����=�N����zhY�5���8�Q��:ϫ�z����1�1wwEa1X�c2��^e�+������[R�����Zf��j�ڽ��kp�vum�k���e���i�c%��fm���6�k��� ��ut�.��eT���oZ���v�V6�7) /$Y�l�ma�hm�r<eq]mU�y��j��� �p��󤓺t����7��fr֚4��������1���^�M���]�쩪�U]4�o�;�씄������$Y�!�桔�{��-�b��e��(2[�KQ�f�Jp�0��@��!��]�x0����,TH��t��c4���7y�%0��V��R���U���}^�)6���w�u�eR9�)GA��a��XZ�M2r��H[h����X��bDv�,8`ⅎ�n�S��auM�,��sD��R���I�6qWVU`�·u�h"W��UŊ�X�,��T�Q�C�0۫�:�&�L��B�\u�9��XB��T���� ��J�rU*�	B����`�q���C}W՛LUs�`�e%!����%f��Ѷk���i3�f��W����U0�E�[����)%n�l�(�u-���O�Ykm���޿C��>I��>sXp��.0W	�(�C�uήp�ݮ)*;��%g0Y�s�FM<3�+���S�+(P�nк��uY�g�YP5��D�t�e�K�Td�F�b2�)��,!��X�*Wsy2�h޺�4�tR[�)�<�N�!c�Q��zΒ(r�sY��OЂ&8!�v%>� ��N&����os�.�X��~R��i�4�uU]n�6a/;��K�˻��*JB��$�D��[}���H�$�� G⒆!��FZ��F�"l.��L\ X��`�A�0�@��ecż{f&��@�@9:v~���F5
1L�Y|��k�����~�ڬ0+���g�)>��{Y}�G[,��t��w��(G����E���û_�		���z~V�BMÀ �4>g��&	��\PD�no���I	k�.6��NrӐuR��GC�x��UT�6����&	Xa�?a�ݡ(�ρ7�~����}�l��eH�L�[]j�R�]-NL2�a�M��0�\�b�5�}}���>��[����W?�vT��A6���1#F�+�Wu���xE ��@� �
�I�Kz�<i�n�� ����`Y_iF�Ou,#��s�D|1/��nTC�X�D46f6��N�um81X����f���+)�@
d}'�)�Uc��N��s5J.���$�ȋ1��yi��d�;	� ��1D:I�v�gY�: ɂ �%�p�*�q׎!��F�X�b2P���#ఽ��S�IN@��h ��u��� T՚��eS��@��%���8a��W#J�W0G�d(jN�I���� �{�m�aCh@Y)88^�N'�̖+��s�0`GV� œ�Z�5B �Wr�q}�uL�%�	"�#�5"�M4��p�`<d[�/B�	 fՉd��t؋����� 		���'̓�zӇ��5Y,I�z����ɥ
�\��X�4��D��O����a۬p~~����eU�on0�i�i)�h��0��C�D}�X��_0�%(@1�(FK�x1���
�����}2���uao��V\@Cp�Ē����T�L%a9�&e3�UG!h���#��7�&�F+i�_̦@��a�(��@�f�\M5�����cm������_���O}i���j�_]9�����h!a�rH�Ӊ�bEh0��of��ƾثP�A�hB����[{���9����/����=imF��eq!��!1�Q1��[n	PZ5T�8`�-��C�:m<��-���A�y�0x�A��{�����4ޢ��-���N!����>|�qZM��\!�0D��*NQd�	t �p���R@=��Tv��&
l�BiJ�}V�.�g�-����ꉋ�yfu�!���eż�*���O��/��1qhn�Ɖ����,��m30�&���R��Yz���bً����[�s���"�ھ����xZ��BDF%r���N�6U���wC��֋��EC+u����I��I���	v�l�w7xx����|"G�k��P@IZW����y�~�v�'�� b!�b8X�1����`@T�)���ϰ�}]m����������A mM�����*CN�� " 0~H���;��� �Q��;S$�g���_��/�;�&wQ:���i�hx�׉;&�C��i��X
E�.� �|E������|(�* h�����Fz�i�]��*j{����~f�$}B��頄~�������-�F_,�����p,������?V����[n��3TRM��wڵ��w\sS�k���M��R���%kْ"�Ў�!��E�^1R@Cj�F�?f`5���ف5F�c������� �W���K�0 ɵ�h?)�in�W��U˖gU2�5���4SBU^���� ��'(@���3��'cQ�3X�BR�H�+b¤s�C#��m�.p�q��M��� �A�|l�qA��.}.�p��H~�*={�����H@���"�D�����#�y���S�`�
(�k|L���n_�4R�����f��؎����#�<ig��j�1�+]h�/���ږ|Ua9�a� 1��6�c�1aU4g�3�'aݨ1��-�ſ*�Ȃ@ė"�0�b9}��������EU=t}��s�۷V��G��^ǎ�Y�U�~��
{��|��b��D2�-eI��=Ci2dN���Y�9u�I�v�]�P��[(@fcg����{�7NB��� YM8<�cG�L{vr�c��f���EY��#�>9�$����:����3����#�(p�a������6n�> l�EU��r��F�W�j�mj�]�*ʳ�ċ�uS>��4{��^fY-w��_��̉��z;��*G�51-�ת�D�@4�e����QA�ڊ�� GՈ�N�	aϊ�f�v�y�R͝�ۭ��R>Cōp�|��<X�)T'�+����BuLq�ǭ`���/T��WR��hR��+�/]t�,іV�&�]p������x�4��z)�[�Ǎ�,�{�dc���	Å�6(	�b���&����[����9s+X���g����������*���S�e>�7��`�qb�q_6�8�>��Wԟk�7|�&ŨB4b�v�M��ˮE�ߝ.-^J	m���z[�ҳ2���i�=�YV2
�Y�c��;��������V�����*dob�P�ջq�p��
�W�I���z\�k�
���7sˉ�<6ŷGMiݮ?,��&{��7�/��|ɻ�՛�aC�Mӷ�.�K���VQNᵛk�xϪ�޳ 6s"�w��V�Ǩ=H�N�4Y��7��)=ț���j)�tj�rrb� �dMe���<���5>~�dX=��e������������T���]�}�x�e��h���];-�|=��Vz
'�3������n��M����3��K�AT�ޕ���r��?=�ϡ�k_h�nfl!m���:���^�r��u1�v/Ԯ�;y3��[�$�5���SN7lJ0��4蜻�x�;��n֎�{�ٝ*r/M�¡�^5	��W���±-JS-٧ FG2�w#�u�~\�-����̒L����k�ɮU���I��'��8e�{�3^����/��W��
j�K)��G��9�c�4�(�n�Yc�Ph:��%���Pen�S(\Ҳس8#��������P����Y
K1�����k,�V�z�ͥf��L�K�����ms�+�7��Qv��4�Lej��Lͮ�AP��ٵ����ChsB��A�Y*z����#�D�LhD,FcG6���(��Ks����\gZT��_WCY�R�F3��S���X�Ը@�^��[�8��(ǽ=~���1�b�k��hoE��?���R�<�,0����Ph��n�u�E Ӏ�i�ѱ�	�i�� OL�.b��++��F�h�vW?Ef�w����ɫ�I��q��(��隒zL���UUM��RTԋ��^2��*k"�Q3P-��g#�P	�(M��z��$Q�#��fc�u�*�{/���r��N��=5b.Xj'g�T�*��}�>{Փ6����Y��2&� �� ��L'U⢯���l"�I�X	=�&�go3xQZ�ꌁ�Ro��p��~����6��V�}H%���7�$0өݺ+������鹎��ֳ�Nseݨ�c�;���~~�\�l���`f{��C�[��TL?:�Ў��a�ٿ�����J�;rݷsoQqW��A��+����}�sg֬K�ޜ����W�k*1��6m�*[k+�%Z�C1�g7LUl :Ì�8J�L=����U�䏧y�x�����٩����1�6��!j���2����=�='�{k� ����'f�u��>�%���,��$'~10,{�"�ט�����z��Z7�n*��^�e����|s�7Q�����uv��Zzg��$�B�4�߫�Y��V�NLz��z��)��,��t1��f��O��H�.��ŗ���[�99~�0���3}�k�U�,�}���ڟ�?���G����߈n%���\Io��&�}��"�t"��(�xF���?�z�R/�^��{J7��v��EϲTi��82f��[�)��K���(1�����(P�)�X)�x�D�#=.�у�Ӓ=fꪝ�����63����`��}��=�~o�=,���g��4
�WU�!�:ŋu�0�M�^P� �҂��*�VV,��3
��lٻj� �Me�:�ʮr�X�a�՞m]u.�os�=+���ey?r��8��oK͘z!Q�N��?h���Uu@�^��֨8�7�H6
Iu$1�k���X#�{�,Gb�q0�ɀ��g.��B� =�������9n��щ_B�۞��}kM:�҈_:�����y7��7���3�j��.�)[������~z���{T�R�t�N�"N]F }ⳮva���ft�e�S�@n��8�;r��8����E�hR�b��W<��tc�M����v.���A9Ld�f.*��f��ݚ:v�m����a�j�a�W<]�)Sl�<��VjY6H;n�;t��*�YM�Y�W�*�w�"檎��9C���{�+��,��v��M�q�2�-���b������ӹ�����ϯn�,A��+������2�^�������`:��?s���Jptù�5eUj�&7�IP�E0��0���p�ޟZ�����s-�^�Uň��{��W�;�~���L��w
ST���9�������b�.���=��!���9/��p�M�QjJiq`,ɫ2CjlS�Ю.#qs�\�U�)ro�3>�+I�yw��+h�,��t���*]�
���fAI�Q����H��GO�B`隫��UQZp mÂ�I�m0Ծ�٥��ǄfTL�cq�=*���R�̣	���]�L?]u���>�f%k�K�B�np�\�|�Tf����O�3{���S�[m,��x���ӞƲ��-53�xԘu�	�<˩�/��*.�-�A��-Y�~�d�Vye�ݭ�z�)y���17�����a9�y|�{O�a!�2�}�"�D�W���y�I
�ts�wԇ�Ξ��Ų�.���.���42�81�W=���NJjc�T��V�u:*��#j<vIHB)�X.�Aڮ�c���B�;��^���˳��.F��z�ߴ�ũy'ug�$�ǻ��>;���|�* _�w*�YSh�,��!ثj'�i�y=�ss�q��,�;#�]/X�fi���l-�e��=IX��enR��F�m9\�Nk�]��=W�#0q���%}�)E�w�V9���E>���I������ �,�-������ߐ��xlﮘÄBV�4;b/�Y������(�?]��}���_�lԜ+���_�P��WMS2����	&M+�|�4@�$��p�4�2�Ӟ���b��B�Vr�ix�q_~����]N�d�|�QN���^�(�(� �Lg�g�v�:�����֛
�b��ѩ��9�x�u�{f����3�/�a[�_
y@�'��U׏zX����K��jlXd����=�)��"
��J�R7&�j�1�ލ�*�_�u�{q�Q�X��g�7�7��Q�r����;N���svh�#��&�W�����oj��H��}��������aI�_�=��߆3�.�3��i��7�⯜c�t�[�̛���tA�uZV��7Վ���ǡ->Y�0Wwo!ԯ��-���EU]�یwh�K�K>6����3T��s8�zJ�NR6�o��jVV.��L{ic�N�םr��4*��	��5��lfYb��˂�gd�MCV���e���.6���M����l�)n�b�t�ݴ����fa�2��6�U�4#,�B�,Ѷw!m��om�ʹ�ڵذ�s.
b��i�A�K��Դ��vK(���7�ҫ���2b��&?���B1�3q�GW]�\.�YKm�8�]t����Ͷ�qP�<�����>}�K�Zy>F�.�ڷǦ������k!Ȩ��|"��E?�=o�$	ed�.<��,���Q0D$�.m��ao;s��E��Y+��l�fz-k����x��LT�ܚ� �+DhM��%ݭ�;�']�ijˋ�v���=貂P�X��y�t|`�C}p�u��{�ѻ;�"<#�s&	MV��ip^��-��t���&���}0�=>�~���l��M6�oֽ(��DÚ^��W�w�T�s:����${�t���P[�.ƚ��+tk<�c�z<50�{�num��2*�zk�iO���9(��,�i��P�
�p�xFM:<��jc~ȟoB>_֞+�G.1��*7�
��@�2}ړk%���AW��͗Q���l8l<�3r��*X2l��PhvR�	�u Q��Ynaa�i�;�����&)��cy��Y�9��<�g����9A�gZ����*�<d)�Y��ݙ�W���8��ЪO����~�U�H@jBN���١�O��ۙS�!qr�ٽX���q)7�S'��$�=�=F�ؖx��@���N{�S<;��C����B�]�^��A�HNL[Γ��u�wQ5ӈ߮���p[��@�p0�o/�QN�],�� �S`�qc�p�=�hP��P^ue���y�݌�|/�A�	h�N�����Ι����m�N��H�N��/R�lwM�'�&Վf٬�Oln��|��mr�{�03Y���s-�5��`����)5P��H��!Y�����7<U�͉	Cn����1y�QM�R5�ɯS���gG�&a�y�����w�==@�QН�==��ϡm��	5Nر�(�b�0M���vu%&�:;m5c��0���\a�~��lc����R�08�\��u�dMV(N�ORS�}�*�8�5�{��M������3x�s�h���I��:���|����.\���b�Gm$[V�����[:�����x��r[���tS����F7ֺ��:6eY���y��(�i4z,�e&�U.�Nw{�3�ߔ&כ���~��������񬩸�F�`�p����m��<��F��ZV��c:�Z��MJր`:�'*a�۹{0:���ij'^�P�f�ފ����Dq:r�ܬKFlm�L)6�]V&����J�~(:�NC�՗ߧe���o���ci̇j����.�?*���A)����r�os׽yO��2�g�h:�4��-��J�La$s��Q7K]q�r�J�cckP�35����n�^!�Ƥ����&�-��^�x�norM%u�j]Z&�#�mV�)�n�mu.i�~{��^��Y�p�� �^=�U�S��"�4���V�ev�U��%�n׭��b��4Ջ�b����˟^�����>����vp���^�����3g�8�fz36�]u{�3w6/��8�� /|je�w>suk�>����j��a��m_�S؞E��k��M��գH���ΐ�7]�s;�יz_v��T�W�=G7ʲ���[-6ZK7���:z�7v�C{�h�����8+��N�s}�m�yc��{��Tm�͘G<��y���6����z�Nm9^��h��K��=o��y��Mؽ�g_G�1޷9I)�pƭ��#���s0�;���^��Ȣ}�{�T��Nto�����B(�'	Ba�;��'�~����*&jWT���Y�92VG���������\%6�ot���]B���@�#$�춓��W	�Q�G�E��(G�du.�$�CKnN�ZB��5�ҷP�5F1[P>&%������M��z�q�{�s;z�F�е1z����3u޾\(=�}��u�fO�)�9���*�M��.	L�0��ⷎ��e���b{jy hT�l���u�*�9� 7H��^>F_���t�}p\������@�lma�Fd�m��LD%����X~��C�[}�p�Kʺ��^��YSe'F���k�!f'��9y��W���h�Y��<��>��Q�*�j��X%�<���$\��Q0� ��Mepl�3A���Qٟ��v��XD�D¾�Y��0Z%D8m�C��U�s�U],y��8f0sk3��3փ��Y{d`��js��n�$�����>�����g�E~V|Ow�n��me�:\�u�r.�N�ɝ�ڲ�Y�nct7Gdi�#�Vv`Ꙏ���D��
S�d�Y34��}/v �����jlǲ��ޛ͑;\m��
�!|��;��J� ���gǨ	W̦$K�CRhA1
RbU	��]L9@����9�ԭ���h+k{Kl�QZ
�WT���L&�b���H0��q�5����jf��&��+�5���-,n�(Z8�HtF�kZ6\X�����n�jk��
cJ��2=�p�V^�[`�<_�>���#4�j@dWGK��%Sie�\��b7���Zw��[�f�[@���W<5$F�~�Y�:�ǽ���D]���)�����z$��b{����~V�R���`x1sp�h(	�Iw��T�/k�]�6{���#����0J������r!9LE���z����,u�ӂ�^�ƕ]���k^�,��C
p������j�ܯT׺��D�N�f�Yܞ���f������
,����|YLd�&�L��M��f��l��h��
L��D�Zh�;�:r��QL�^�\�\��7��Y�~�Eh�^�E�T�n.ѐg0�;�0֖����|$I��@��-J��ɘ��.�0	�L�*��<ө�����P���$o_	��遨8��`[�8��y'd�oeׯ2���@ey����fo�v=�ϖz�{׸�݆V�0�깉Ԅ�&d`��6ˎl uʔ
3~>>��P�����|���r��NvݡO'L��[�Y�:�+����p��ǒ��Tit���V��v+�l�Z$��^��< ��1Τ!�O*��]��Uc��ta5���9������j��=�w"�5�x���QobM�W��Q��l���i(8pÂ�M�1�w���~ł��k��-���ݯ	�xB���s%��|!�<��w_*�s]����b 	�%�΍�=�y�p'�\2!$�;�|�"b��WO'��\گ��'8�N�W��:~����+s��|oq[:+b����}������T��np�+�"�;�3X"n�&��cX�?u_Ol�ϖ�T����h���3Vv#���!:�(����ŀ���=>����jJ-:���@��:l0سm�suKKYu%�c]��h�R@2�`��=�bvx%�Y�t&H�]�NC�P����|�E,��q�t��`i�Y�&�օ�x�rS�U��%ӽ]pd��:IL�m2�Y�X!�듑rX;$�+T��.y���Z���n�tͭ�2���\�ͨ7������q�,������)^�{��+ߏ��u�;��sڍS�>͹�°:K�\�nx�]ޗޝթ-+��K[}[��b�o�����٦�Nd��݆��؛��pt'��|�(6�7L�r��9Zq[��X��Zȳk]�-*l6݉���+z[�yV���3���zf�u�W]9�kB;���гJ�#T�U���5�'s�hl2���;W㬘��{L6��{��TqW2|U��d*E�{^�<o�ז��=f�S��n�R�W<�	�U���u�_��HS��m&hnC������ݼ�G6�����񊮸�ύ�w3�o� ��:����4��^=�$�nǠ�Z���A]M؇#���*p�
��`�ŷ6��u��K)3�E�:��V�r
ܛ'����|��ߞ>�}]�6p|�70-ŹGm��k����8NZ�Zo�����}����x!�S�fL�UD��fW�Ӑ�.[��g��ɣ���{}q����h�F��[�j���)��K�D����s���}�k/�0E��Ԝ�!CA�	E#֫ig"��W}�R����l�T�Sݖ2�
:�]�r��zzMĺ������{ts�P>B�ɞ.{���N0$��Jw�2��յ����S��X�E��
�i����(��th�j_O>��mL�T�x�|�z��;Z��f`��+kT�[�+�h䙩9�(�,޶�krc-/o���I|����F,��uމ��	�ñ+�aQ�V'��e�6�Ku�blir���ȴ��F�ٔc�ۓ,f��b���W{�)Y�^��mn��5X�)Ļ�9���ybصY=D�D�r�P{�8{X�f����Qnd븪ުwt��RÅ
jP�RN�^n�UZ�|]m9ٍ�n儻����S��	J45�*�Hn;P�Qc��ЍXf�����������g��m�����[��T����:���\i�	pxg���M�,�˪�7��!e�KƎB�!HYV�W)�T�/:Dj�s���IP�	B*�
G�Q-���V�e�1�Si�����τ����̖�R��H���z�ov6�\n^�_:�tL�t��)6��ڵlrpn`K�U������R��9j3�-��|f�µq���9���9�J �<b�f�sס�M@�	����)%�@:5@�`Sr���7��xξ�9�+�f�fn��(�s)�ZS��v6���D�}��dε$\���Ζ�FP��R��e[����X�Me�$��
�c��Gd[�[�w�i�y7ך���̦B8r��#��m0�f�\4V:��l;r뜵��qGV����M	Kk��h�M�d��rb�B�ؚƃ��Z�o� B�R�;F�Qfw��[[cb��Me��ju��K+4).�!���]m;=`�v�G4�.���`��/ΉX���z�~o{߳޹�(���rj-.� �ha�mG]�Ësc�P�t#ib������I@b����"�3j���8|:-+��v�8H��%�� =~F���Y��Y�Q}
_�\9R�0=���N��k�ڹ�;���������6d{b�����Og��e��:��ʓAo��.)f��9Ԫ������6^��-4�e��������3}3�S�q��ހ���a���q�1�!�*v��+�VH��R���%;0{`rJ��	8`�Y���s�L�f*�Nf�=��n]�
���>x��6��z*��:3콙뻃H������nޜ{L�MZ� Z�_��$�E]�I�X�U��O*��w��ͅQ]GK�0���uۊ�5mXƈ�[36:��X%c�&�6���P�F �9Oͦ�f��dj�ջ1��Er�l�����234Ŧ&s-���sOpg}!X2��)��h��ӎm�'y�EM�A:6bl�����Ě�n2Ը����!Ym0��z��7����O����+-�����Rkmf�sw3@��\v�2��4��h�I��9����J`t4����E3%����A�u��l]WR���n6���҇O������N��ރd{�U������z�Mu�@ӃȆN���Xo���);%�{/�C��ך��=ю���^���n�M96���p/�n�/bX��{���6�v7[�����%��%���*&'�bd	wJ�j�+:���:z�0վ�����W.�dWu�����e�'r\��*W*��/�펌�0]�M���mYmka���j�i�� \SA&�jM�f.���"j�J�қ�T������<��;����ch���X{&eh�ڲF�Ci��/"�a�������'\���-뮱��tw��2��o���+���N�n0k3���Gܠ<�r夂���x
�7E%R�eFe���U�J���}L�4tv��Q�����r��<}lߖT�8�ʈ�b��4^��)^� k�Y�e�s5�ܴ�F*��c�q��a?�؃FVس
�tڣ�����B�r�Pץ��fQ*	����݉�7�m��uަ�1-�M�]��,�x	^=,P�����^Q9p9Ă_P�E1 �M�v�v�L��p�����x��xBK�{g�Ɓ[���Sû�'J��y�������4��q*�ӿsH�@80�I�p(闦	�yV.�>�UN��EB(�z��LC}�w�xum%��@��=Ԑ}wd�l��*�$FdwR�=�>���m�������m��ؔb�p�1����`.��ݙ���+����e~��oߞ�����~���x��G��\��$�kf�������2�=�J�{�L��#!^{}բ��p�iʽ,g�����qw0��sX��s�>y�%�}`�m�j����,R��-֩�*զ�^�^�jܢ+Հ��L��)��M��vv�ꢦ���»FN�̝�l\R=ť��}8�{��ǒGK�����>����i��ǁk{.y�*�-�7x%�U4},;�����+�@8eQr��6������o�7��2���T�N�7��D�AJ1Mɬ\��P�L�kl]������rM�K9-�����<��7�mv���*���j��]�'��.v�������O?w�� P
j8!���j����24�3���l涚6����K��i�d�6(�+�7�ʊtO<�g��_}:}��_�;�g@�/&X���a�����n̜�̇2f5JN�3��e����j�A�}0���Rb_1���-	b�(��b�'{��������GU����1�v��~5ڕ��G�.�fz�(_2� �sT%�d����.I�׮�'�L��1�"������n�=t����K�^᝹b�>���|#��js"c�U]f����-��"�,m���X�l���J�M>��@�"=-�]�j��wu=�8���Dˆz	��XǛ"%��en��D��(pa���ː���~�����^�Q�eg���V�� �"^�_OH����O�L9��<5����?����H��/�UX$�	�D(�q:�Z)�<u��*i��UPD*Ie��z�8K�X�$8`p�
"�L�'��C�!wD��T��THP�����i$ O�a B���$��I-����p;�L2�����k��o��d6n��5�<��,HOg�s^?u}.�Ӎuo��Q��s�!���Sj��Y�?
��~�5{x��
�U�wi���=��C�io��m���U�2��ð����#�����-�s�w��O�u�����oۢn��9n��x.�D<�,
� �P>2�"O�%���wv��S�R�L�jL@�ec���O�Lz�>���>�0�}We}�k�~�k��H�O�?����L��^��0��>�O��Pu	t{U8���'��z�����z�f�x��<�����s~�`M%At_��O�p9�HB�B�H��HE�!�� ��B���0�`*:���(��%��a����BD�C4*�j�0�����S7唦W�20t^�L=����u��ɒ�9lɀ�m��
��%u2gjm������vfg���ᖲ�"�|�XA��0�0o�A<6s��ڍh�(b�sC�D���9s�G
����F�,��xA��D�C�PP��>��RL�����5w1�T4P��&� H@�į2�0��w������� Q=�ۖd�g�,��4�ǫ*��B�qP�,��3f����4&�U��M��jI �*����������P�B@$��Bv�5!C�����_�����1��1;z������P��@��
���ϳ��F >���O�%�"|T��5	 �*~����9p3t`\U�i�J�9�R��	l�a��F��Iot�~c���hp3��{;��fN9��`��3��X�l4��s8�$@��#�zL�|6�I�����]��ݹ;���}�g����
��&9��Q�0C:��Fw��S�-��o����֠(�1��*��A���}Ǫq�{^�?���>r�C�$�vN���]��BC���