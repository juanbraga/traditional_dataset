BZh91AY&SYco�� 3_�Px����߰����P�=ӹi���I#$MM���@i�h4i�A*i4���A�# h@0�	�OPh�&Ѥi�d  24��A�ɓ&F�L�LH� Sʞ�<SѤ��y@   �E���"H/O��/��W4P�k����Y�6�V������{�VU�J��!�$E�ݹ�aͶ9���շV?�ƒ5<Y%��y�,q�G���lh�P3T�@J�	I(��8.���s����Wh���LY~X����,�L@w/�o�l((L���u��,�â�vA��J�y������`�y���t@���f�s��66���� �;���J2�����72�%�gl�}��	?СO�ę�%����Q�5�V�:�xh����x�5I;
�V��=�忰���?�o���uC>�7
�S�a��ʥqr|-.��7����܀�*�?v3��cy8|���ȲH�ͣ�F�T3�3$寤R���b&���ZtD.�#�<%����_ݧ�X�F9�KX��p&���BRa��ӯ6�gn\AaJ7��1�a�i٩]M2,��G����@&OpM5Xɝs59#Y��L�4�F'mX�C�*���[��5�D�Mq ����$}\�����b8ӗ�%�E&L�juK�K��NG�r�A�^a0hk�H�b��8��T��J�R*���a4�4��#��D�
ͬ����w[�P�[%������j%J�"��$��N��JL��'	��[�A�hU{�ʧJ�"��j��X!PB��n}�zM�΢"购��-"�+����LS���y���3���q��* ����ܘ�:��ې��H�r��< �G1��B�"�!��Vd�&s�2o�em�F���q�E�$�d����NQ$q�E�j�EL)A�$=���
5�r�	���-;
�Z�� Z�CJ��R�X9
'r�~Ve�^O���n�8�&A�knX�rE8P�co��