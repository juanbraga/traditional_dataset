BZh91AY&SYT�֏ �߀Py���������P�m�=��!J�قI D����j   h  %	��"@4 ���@ $D!OJ0�)�4�����h��L�i�����a�0  � �a)�y=)�h�SL� ����13�UbD�Ar:�'2�@~u%�f��Hu��p4B[ �G��r�Y��t������e����3��SMҝ�5ⴌ�
XM����Mǈ�ƶʘ�?�d�����I'+� (����b�*Ud4��c�o�z'�d��2ftv)	]r��ٟ����/;���gE���|t�X�'�b0��k����G��d�s���K��-K1t�]^MS�d�][��U�'��dŅm$��V�+'#����5�I3������-�����l!��u_�O�E�����M�G��f�2�&b�t� �u抎Z�X�� ���@ô�z�$�6R�\،�\�+E��֭�2UR�3ry�Z'%�y{q{4{{�c*3'+��C:*d6d"���b$ϩo��ChTQ�m�=�Kz(��b[ӳ�Va-f�u�P�5��j�E�f3m"�r'
�`(/�9.�yR��c��$-Ns���T�'m\�Z�g]�cHª6/�$ݦ��s�iZ4M#jl�Lr�,� e@�Q
0��50�Ѹ��� g�P��\Ù�ILa�<�>q����q�5P\�
�oYk�%�a��N6� ��us�I�*�=+�S�����S������m<Fg���Gŭ�q��X~o���A�m���x���k\��N�%� �r��őA��(�I�Y�,GaD�n)��p�k�T�E$�2+g �/)�E'%\��τ([�A�b�Vn*ZU�6�2��HH(.��ѬCl�A�)�!1iVT+�G�%������1�Zp��qfH���dw�N	Nmt�D1��Krb�Y��2t��OZYN�p��[c�H�e���e8�9�+�#�H-����c��Ik�\��'��"�GX�Q�uPPR3X�H"��(b�����N1qB���U���^k"B�E��V'vH"v}[�D^�q+�Q��-�$TC��_f]E�I�व�j2dO����w$S�	L�h�