BZh91AY&SY^۫� �_�Px���������P=��.��� �)��M&�Se�Ќ���4 L�@��M0� �� $"�I�Sʞ)�����4��4Ph=O���b�LFCC �#	$	L��������� � ��>��2hE$� ��(��N��u��ďfmx�wX�i��>�[�����q�vj��Γ�s����F�O��gn٩�Ǘ��dA����Pt�����˒.��7�,�k����kq;�О;�f�j��@)F��8]|-��g��,!�&k�ؿ��$?��|�	��o�`ɞ�]��<·�G���GE*����(�Rt0`X�D'0Jd2�FD%vY��{��q���Z;U���1�1D�X0�n.����E�����aYL�{fͤ%9���3ek�l۴��&�c �2(��߂2\���Eb/2Tj��wx7:<��zS4�6l�[\%�Z�*k�F$��-�X�L�%��a+���w��nm�����4�82���������qe`�V�u�_F	Xl��YVtȡ��X��m,����5A��ӏ-�̚�(�36�,��v�[Q�Jz��`����������=������wXRU*2ۯ�Z�m�������?�Ż.��5T9����lm<�%g��;�HG��;���o�wmc���B�3Gx�uo0�8�g�2 �q���|>��3�����s�������1(B;"Կ��b��L,L8+��.b�`s���#�WW@!LIs�p�������F4f	�O��0_(�I�ȯz�,���J<�%d~�q0 g�Ӭ'��)�0y�
��x�&����kLB�iL�<B#�釬I��>�D�,���p94�Vi/�ӉYkޜj���Ѱ�B-Uٙ0�&�#�����4c���Xp��lD#��<�k�a9�r�R����KZ-^��A�+"�HE��3�҆3ߐ����"��K�Y�n�]&U����F�Hr �1m4�mJd`�B1��rԠ�caV��ÒU�V�\8Sk���3坒b��II�0�5Xqh����8�:�w��Up��Q✵A�U!��"1D�Pk�f]ND��f$� NPR-*�F��c@N�S[)DB(*Mzk�ZZ�8TŅ
�%"�0�5@�=������b�1�0e-���+;������e�iQ�R�_a���6�d�t��5f���"�(H/m�� 