BZh91AY&SYX� �_�Px����߰����Pqn�#:�i40	$��F�4h�&����4�hh�d�~@�J����2d�4  ��i4&� D�A��  ��A�ɓ&F�L�L(�)��h�L��I���=  FL�(��Р��PBE[�F:��ڊ�V�N�R���`G]EDl	��t�����>�.��F�@���I�}�-��8�91��b�Z+���ձ��T�J�r(�N�駜�5bƛn.�l�CϨ�e�ږr��Z���
��p5[��t�H��hؿ�����q�Q|�����`�����(�u�g��ZI��!���Ľ��.��H:ì�DdqdA'�xe� Ż�TP��w	�}bd��q��@�)�x4�Vq�23�hʳ��#K5gG��JA���k����:��楔���k.�$d�`�mfb,䌜K��)\d��GKS���ɦPt�kjn���K�-�)���p�$	|��i$82��x
�M�V��\�e>��f��B�m��CA�k����#ƙE�!!��`�xg�v`���n��0���8;���MO��k�цn��2�Oo���N��ʜy5l��P��;��s�$��n���<jiq���4L��r�r���I�>�%��]]Pw�5�"N�3!��(�r����"	Q�u
7��������
�Ǹ��8LFH.)�}��3&h�;�tQ�h���]1�+�W!��qr��pj�y͞zm�`�\`��#%�����gGpȰ��d$3����t%��r�m[�"�t)�Wc�4�4)��6�		0��e��������)ӊ����u�/4�_�������$4e��-U���0ΖA��?�Ȏv�Yg����)*�h6�<G�2H�.9y��&
�GU$7ʷծP�I
XT��!��ͨ�\����l��g�)���\��rV��-�Ci�,EIJ�Kq�]� �;���M�hj�l2-}Vc7x�����2�	�&}�H��r�����̶�#6}@`AH�Y�gw�\���km-1\e<6��Lm`�9V�ƌHA==�L��aFZ�*i`Sa@:X�RL��"k}&�*%V2�H�!!�3^�{ɖ��Y8+be*�e#&����]���26�,�Ț��Ǩ`�-�nU+��2���If\�u
s���6�\l�,nV��O�.�p� �)�