BZh91AY&SY�9�  ;_�Px����߰����P^\�����jRD�4�dd� Eʛi�4~�4f��S�'�2� i� F LLL �$A�z���  = sbh0�2d��`�i���!�E'����҇�(�M6�C@ @i�4Q�R�tQDID
�~ϓ� ���)��-��X������drd�,I�����܅��T�
)8���%��<+/e�!-i��6i9{:b���;�4ҩ�<�p�č�7&q[���%E�y�aCd��(юb������8�		�dϝ{0�cg�a��tdlѿN�|T�8Wr��� �Oo4�m�ta�iY�"2�h�BFP.�^�� Yde�WDj�% ���Ӌ�|�M���drj&B���S�E��4��$�*E�d� 2�G���l��g��P�E��%��b������1H�ʋ�,Ů�Bע%�l�$DԇHpD�J��JbnhJ�/p���������,�M��؁��UNjeJVx�jݯh줂A%�I � ��sw�9 ��",(8�sBWv�"��� '����e��D��� F�� y�)���#dc̻`�%s}�bo��^d�����9G����G���������c,)>5�_�OAP�v�W��^,���������|�u��g���AȬ��I�$/��n�d�ڼ�۾�3[$@��1	.�@���-&�R���M���lg��H5��z��0~6�/3APiqQi��0�d�ay#��nP�Y�s�Tb�7C��wk�����r��P� eaa�(3����4;���hE��j��IH<�u��r�4���5�ӄ���1��ܶi^�GySy�B�S��-��e���Xha���O�/�� x�j,/+�_�D�Z�S�;c��:m;�B��̘lu�6L��p�����V��+�Q��a+���JAP� ��L%�k�U$�
\QU��"����Ud���J�C�����:
�t- !Xg؍���T ����6�#�۱��(�y���f{h�Om!��)���c+��~��`�2Ln7�Yp��`�Fx4�"
D���$Q�m�Ds��(�Ni�uD�DXb�6�x�hP�֟��42W��Y���^��I��Q
m��E�
H\a�.ko���11L�H_����e�띚_�e�C���}Ljً�`ِ������\�Ӄ���
ֹ��fT��a��ӽ�J!�ח�k���H�
g=� 