BZh91AY&SYe/�e a_�Px����߰����`=��M  �e���$���55=2�5= �L���� 5<�)ACA���     s F	�0M`�L$ԓDiF��A�Ph4   s F	�0M`�L"��Sd��y1&��dڀ@�h��PC��!�*2 %�(J1����SU� S�.����$�P3LQa�L2b����>.f�41ƚ�5k=�\�x.�'��~?��x�gUSq��,�;�vg�;9wdX; Y�fdJ��Ad��#�K�����nGqeL��]��.���S��0Z{�N/�v�n!�S[M(���	�`��4+V�2��;Жk��&\���8Te��_��w�A��w��霫���68�JSѽ)�k� AL��H�|:�>��؎�#�g�{�1e�bq��s�ՓYUY5�wU�Y�������C��<� �Lڟ�6��m��~ǻMե��~��NX��:�RO�+ʹ4A%T̰��	f���	$��|,mi�p���ȡ!\OE�P��N.\��*̰�1dԺꕆbG �9DL��q;+��ج�1m��8v�8j�q�q�Z��`����T�"�ֹO=.��[��u� �,©\JaF�ڈ�F��Ʌ:��ֳV:��v�"$�mᙸ�d�̽�k�r�[��M��XH��6~�ܭ�U1(ɉB��������[��K�5�*wm�-l9�[Ky7ӿE�@�I�����$�uyTn�&�b��rM�������3sb����]6$�8�a�$I$��&�KVa��m�Ȣ�Zo�2�w֗�SzB�689rM�{i�Kܠ�Y�]�Cj"�<�����XЙ����ũ��a���V�%�jkqQ"�w-L��[2�֧ݭ��`��B1�补Ĝ��y��ꎆ�ʢ�<.��k$���S]I$�5tƣ��K���".,ӵƬj��=U��JKH�tE<�\�-SM�;fÓ��*ѓ*�4M<����pA:s)�E�R-9���4TQ^%A�@hK~4�-�i;�t��,�u�P1$1!����6b��$��0PX��e�0L�d,Е$:�B �Q�S
��e�Аg�1�7΍ivb��7��Hh�8��u�w[U�F�K���=+���o����J���ǻ=��bT�����+nD\;n���Ш��T�*�u``D����: 1�0�q9T�qol����krD !�1	.��l�9��)U���8rHTw������i C�������E�`�(b���&C�j�ὦ���"�'J�m|�ǘ���1�j��pc07s�s���@�^�X0�c4�B���Y�Ì�)D� 3���iF��*WZM�S��h���t�#	]��7�K2�q0�] ��YF
9�k�]�ʵ���,���XR�\���-9�d݂pҝ�Qi�H��fd�h�?��^m)�+�Y���t�#@]��1��-9�5,x��$/*�^�U$�e,*U	F]�&D�a%䥣Q=u*p�M��ɫ��%�d)l�N��U%j�K�4y.-� ��Sahi��/_E1��C~��&�8�ͷ��V�X5͙q@�X ˛J��)j9���@��M�K�qZbN��ST���6Wi(���h=:�_}yk1*Q��>���ZJ���T�
�h  ����M�l L�&��&-0"�EWYv8�+ >�)����/G�Mgq�0q�)V�b��L�����6e�`��gf6�-̙-���lZg�rE8P�e/�e