BZh91AY&SYs�#* �߀px����߰����P�8� ��	JxI �4ѣH�&��S���~��4�C4���AE        �~EOT�=&��4hd     9�#� �&���0F&$i�G�A���jz� 444ڂ�)��DS0R� (;UR���������Z.b�!Q���>ۊ��+�H�x^Z�m�������:���G��ig�s��)��\פ�Gj�&(C����4a�	�D�L��� �$�6�K��o�yD]C$�c�ϴ��+o[ �:�@�N~����rXuO�@�g��{<�b"�&l����F��u75%Aq`�|_��sNyh��{/
5���������f�8+Tms�;� �8�Pg��H�����N-�/��
˹u�3���a9E��̘��ʑ�b�$Ԩ��R�"��@�U3/��˄Bp��d_*���riŵ8Y�,�J*�P�uI��.��H�i���R`�)8cl��[N*�mC:y��v��ͻ	��F��4���P5e�D��ND,�C��e��k�9LEC�ڹ��h�2����m]���:#`۞}7 �V��x�L:��N�N�՝k,���.�{��i�HHI;� AD�B�޿o���r�-4��+�􀮶F�
W�Z���M,b%V�D������FRe6R�3����1�O����T쳻?z���{�����<�f5S.��SR��V���ۄ�T�??�?8̈ԣ���GX�E���I�X���S]�o�u=H�0�
X�d!!ل����U��u�DR�)���z�r�2B�x!��ެyw�-41P�p#�{��a�a����l�����aI=�R�S��s_�J�:���~�)�~Qr*=$D��).S},n���Am��7"�(B�T[a.���I��-Oz����y@��DM��!������06�l���Ĳ���5p��M�-R ZC����iDڹ�b�ȑ�k�Zq��Z��1�BY{3&=\�9�{�J��cG���A��Ԫ��"'q�>4֗�����4g3���Q���o�J'1m�0 4O��m^��Q��e0�)�ps��X3f�Alգ���(�����n����jB�Ga1s�t��\[�0����W�w9���`�W�o8�r��xDD��z���Ҟa��
DJy�΢4,��n����j��L2��s`FH�TZ��_^�S[�KHն*�b�����tP&�WkE3n$���������Sc�Q�M�]�Ć��+C#|@�iFe��4.#wM���V�is������{M�����l[&~o���"�(H9�� 