BZh91AY&SYb�y _�Px����߰����P9^n�r�T�J�$���=�OD3S�mC��i�� h5O�Bb��       &��y z�z�Q�@4 h���0&&�	�&L�&	����Sa=$�	��444@4��D!i줅v�D�AB Ȅ�	�Ϳ5�.n,�&e�C�gF�KHİ�dt1#=���f\:�F���e���������]�A���$��kc�݋��tʇPwh�b�	�����A!��*�gΕ��L*h�BX6��.��5qZ�	��g^�����X�ZL�I�;{,ֽ��6|�,��{�Ќ'��J���n��3B}�VxN� �Vn7vNٻ���Q�P6��/Tэ���pE���'N٦Ĵ����eZp���.kI H{�w�mS�OL1�D"ىJ��0mh)��V̮m�ʆw�4vgu4Q%�L��0�����p��c�ƴ�X'�;���D9�ͳ�������cco�� N�NNd߂վX�/5�������+�L�f2���]���4vf�9����Mq�5.��c�
��1T����-?�����2��ů��o��������Bc��3��g�����ޚ�H�͟����c(��n�����f:��0H����s֥�����%�N�6 ]�
�H�/6�=�N(�[�n�	�q=��f�]�B�l�]%��2�Ir���
q���%�'��{�DD$N�y�|m�aW?w���:��{ݛ���"V�2�J�!��XD�G!aqC�@�X�d���ҫߥ�.5�(��$�� P%ڴ`w8���L��BE
$�b�:�iȫ?3G����v�R���r�"��)�[�S��r�yb���@�Q.fi�,r�w�(":eET]
�P��B��6�������&�P�!�$�f��M;�\�	0�o8�zE��TgF�
N�>T�V�n˫���eA�[2�d�H�2f:��|*1�@��b�׼`���y>���}�h�8$)��&�`حd��k7r�L��r�c$��3,Cd.Z(:�WVOɜ5�q�F'%�"lk�F���hDSRx�p2��s���O��)�"����-Sd�p�>R52�MBK'p�C�300EM@Z�ʕ�\S��j�}�@�p�J���`�Z#��0`�5�ܢ�r+2\�ND�E�v��g��>��ld��d��Y��_�]��BA�Ƒ�