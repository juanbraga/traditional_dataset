BZh91AY&SYc��� (߀Py����߰����`_�ݏ@ ��D���� �'��LQ���1  Sd�H4 h4    �{�T�M�h2i���@h� ��(�@  �   h��2b10d�2 h�00	��oI��'��5=�z���m'�N*��8��@KB(� PAxy���������5�x�����KG��tiK/}y��8��۩JEY H �`&�DD�%9�0��HI9L�I"�2���L�?���Qm鿭nxe�z�ل�o��1��ql�-�)IH�=���wfd'�蹢S�A�E���I�K*�es5X�D�J3T'�"��10\��!�<�� ��b]L8�R���}R�m�D�`,y����=+��ww����_{33/ffff^6>ffFfb�˸�j�������9����owwoy����wb�332�e��]��C��<��TTUɼ�v������+9�3i��������SJ�J{�A^E
 �:6u�$�I�%����������&�f\�]��:.L65:���KcFd]�n�s�ou��8Xrz�K1'g O:n�\v�b6d�ƵjXm��	�/�H`!��oa�ru�����=I$͍ �ċ������a�X�*-��&���;dv0����4$���s��s��$�IC��z5p��5�0j^C\�te�X�rWMQ�k�@C� X���m�`�rI$�m�@c0�0q]!L�p�>�.��1��L
��˅�9K��1����G.�7Z��d�$�pݐ�KCI��R�6!��n���|mCe	g��{Of���B� �I��$�I����T�ȥ��\���-k���hwR��J�*1��L��$�I,͆ٝ�f�A�Q���Yb�5��*�����,��ki��F�=�Q�$�I%\���t�� �WQk\>F�eO�b�*Z%�,19�'�"R��RIS�M�����i\��ۛ��^��.Z-ݚ�*�J��,��B����4�W%Ph@W�o9M���$���+Ie_\��ȅ�Ő�(6�PT ���


���D�
���
� �HJ"

�� ���V�v$A,@, ��M c鋖((�Ud�_a�< b@e~�qZ<?�ww���sW1�^ϫ���߇e���:�;\r M*��\�r=���~5���>xt|t^b&vQ�4���)^۟뭜
r��r!�@P�!|���u`������S�"�t@T_"�u���@��� �ܸ���L��=2P\�w�H��3�xnw5�!z��7�,�nln��.\H3��(���y�k:��i%��hTj�(z/ �#����B�!��.`��aһ����ى
�.�2'�n���f���tP�n��jmF#e�O�-Z�8��4`~mͣaC#7&\�̪ͅ0[.~��iPDf*��-��"�N���ki9�1���5�� ��=��a'_b�dO����5��P�2Y[0Y<�2),Y	�B�q���U(&��'	��(�d�Qr���Ы���T
�j㼰�Pw��ڀz�$��P:F17��;����7��rX�	��<5
�ʘ*L�n;3�4c ���p�86f��6� ]5�I��l�$���U�HXf�j-Tk��iӤ�p��JR�h4-NH��r��8�D�)tW E@\K��rY���B�\=/�p)�D�c��ca0T6���3��2����!B�0�����d����ʆ�Dڨ��?L���H�
t��@