BZh91AY&SY���;'�_�py����߰����`�R��          ���   �    � � �S�    ݼ  �� (>��"��{n�5�tU���{2;��^��p5�v� x8]UW���e��H�Z��d
�����g�@�4a�@����\$uP<�GZ��F��Ca�� \  �AOM�p�h��
��`+�r:�7p�P((;���h��  <�.

����h4øPH�05�6=�A�GAAr`���h �� ������ �h�)���B�AA��|�P (  �y��*��&ML���@dO�4�(L 0  �~5@*���L2#�0!�Ob��5U4�     &�I����@@0�� �$24'���OM'�46�M��v�!����8]{lu�*�a��u��m�7�
��� ��OԂ��D�~/��s����"��TA
�����I��H@؄�HJ���`�TE�.Q�n�㰷/?7���CH )	��H
HAI
�P��KAP3��TZ���H@4����T M$�BEB)�"�I R@!	1 $� ��HP �	d+��f��SAt�ف/Nv~	�O�O�{�?3��7��_��E�3�Pd������ز�fV�r�Ͼ�V��pPw�;~|�#Z/R \�J��Ys�
��R�u�}�ǰ�5d0Niv��:f��@�����q=ڳ�����"j��Ǥ�s�Wl����WO�]��?U��)�Y�W��7s�l5sΊf�=	]t����J{{�ѥ�T��wVֳu�;w:����<�MUaK[�ȓyV�Yd\;�6���^2� �wt�{�`9m��l�A�2՜j%�I�c�rƶW��O���8�����:���fp�2.�u
������O���$ �8\��B �|�3����3�s"x�X�(e��N�0.U�I�BZΊ��s;�G�&�-Fl��B�s�\�}T�o^�|�)�rpË�Sȧ�]��o<��s����Sm��@���n�3�mu�Z� BG\���;h
��{����w���%����;���Ǒ�u�waa�m��\[�!�"�k�u#�`u��Pp��ے������=����{���󜓲��a���zG���Wew��Smc���:�
-T3��Sܭ�S}v���a���+X2��kႫ8sƝ(���;�`Ʃ憁�[�.�T(1���Z����y��jwF��cx}c�{�PI�����ر�\Vi�ש
������F�5����b�9WF=�������:hǔt�6( �F���u/z͜�*)p�{�'f�IE�Qݝ�3���;-�[k�dnN]z�U��Q׋�ކ����+��Ա�^�����9�ˇ�J���.:4>��]���d�Zڲ����\EM�bͅ'�eg�O0���pl@�MI.�����-�z�;�ܵ4��ٕ��t��1܍<�!^G[�\Nd��+���H�>X=��eXB�v[��*�*.qX��ك��к�N<莛6Γ����v����'��Z�p*���.43�qA�r*9oQ;�{�HoE�؆hLtz��(=~�ܱ�u#o,�ћ����c;�K��;r��q���;i㰂�(=��h�=I��i��&����Q6��/ǉD��ƾ���԰���g'.�/(�����:<�*���Z��������a\��ȞC�ԴB��a�cE�'kĕHH��QI�Ϸ::(���Q����5Μi�3��]nY��{[���e��wnP��� ��Ӛ.l�]y1�N=�{(�B�홹�q,j��W'm�㉞�"��l	مVkw  ��sO�t�"ȵ��K�K�ӏ�gV�X��+��i vޜ�B��P&n���݀�pb�F"P��-�Q�ɬ13��@��F��	%ss�J�O�op!b�p�.f�Y����7�˳B��ņ�ij)J������_f�bOh�����ާ%�ͣ�Ń�f#.�}W\è�"t8�?�ö9%)Gj��*���6��)C����$�y3�kq�⺇;v���7G؞��o�����,��Nޗ���Ύ�p�H�^���O�nk�*vm��,}�� �dh�l붽N#�p��Wn9����c��r'���pb�h����[F,����@e�|�HJO;�L�r��S̝N�ɏ�v*�u�P��9�GoO��֫��۸p��GmH��sGqW<�v.˼���\�y0���`	�����:Wv�m���l�t��s�L �1�+�=��;7�%�$Y �'׀�&��q�:����n�Uۀ�"pn�:�M���F�����
r9w@�7�!�u�; �g�}7{�����ZƊzP�t<jM �p(�noo���`װ�gu�;��p}s�2,]�k�\ͮ>|���8��Lr'{��.��;���q�ȑ�p�ԺX��w����ȉ�sR��j��z./����ݨ[~��WԠ�WnU��.(O]���(�� �y�:]�f�	�wT�]�:��Y��,�qó�P6�R��bx�����8��`d�.J�ˊ0�[b�"ܓi���霁���T��9�v]��4d��X�f��]���hw�N�+����c�k�.�
�"��/�@H#�SL2�$.���;��5���і۱0drka+����������*_�����}�Z�ڍ�h�Ն����WC�a�@�]��t�W<�s��ckz%xC�(/��z���*��,��{�f�]����;���kvy�v+��燉��N��^�Ֆm$�^�������&�'��:U��<�Z�˞��+��޲�[��������3�d�y�^�Z=����>-����˺�eȗU�]L�����8��R��)�=�5�Nv۪p5��V���p���]�֟K�6��8���8w�S4vu���~E�8�u������Dh��a֨W`AQ�:�|�6�5�x��kfA�M�#n� rvwff���v,t��I���p<,�A9�\�-�mi�g�m��m�;i�V{s����������=����[���u�����1��Ը���\DۅX{p��nr�p;����<ON��Ħ�o#�a��9e[\���W4j��=��p�\ۘK��*5�cGg��Zgz�pVf!�7:��===��>�P^�b�B��.�4t��	�n�N�Q�"vɻ ΟN��d:-����s�W;.�V�8nۙ&��K�W�[1Fϵni�-�4�m*���`�"dB��	��3�P�M��j�X�!�۟nx�v^�3R� lj�).2�P��z�ǧ����vy�t6���o	�1�<V]�5ҋ�K���u)q��	�Z��籀��n�����xl��z2l�[iQ��d{uvݲ�g�,rl��c���F�[{n��N<�ne�]Tn�*�ku]��RM��[g9�+d�]��0&ݭ+��+�r�rA>�Y1ǁ�P�4Zݹ�`ʘ���U���8$y�vɳúŏ�	�;[�}q��=�F� ���8��Ss#�]7O.2-b�7����xCq�;�{M;n�	�K� �`�z�{q��6�i�є{{���-�����оL�{6;�Y���vu֧2���c<��I�ς-��ۛ�@��H�;R��F�8��6���Ԃ����9AS�woс��{m������뱳���:m�n(�AD^M���=�`�B�qm�n�v;�.�n�k;y�H��#݋u���o����|.�vկ\�{c=�I�<�ۓ���g$��z���n���	��؜��h�'t��^L��q�xn*���`��[I�[Y:��k��m�݉z���=�[:[ga:��.�=I��4�o3��v�!��Ě���^�ix�8�xuѮG�mU��y\�{�U�ӱ��Lan�㌲F|�n���C�nzxh:立��lt�g�s�g�7;p�Tkr�q�lʖ��MɊ��ܯ;�ֶ�+�[�k���{;��=;V��'=\[=�[��.3sې�l���v�q�]�<n����9���L��� m���	�R�xc^���ukcx�n�m�p����癹��j�n���ռ���/����g-�v�S,nN1��K�9(ӽu�"���G�_���)��#vϓ�qɇ`f��u��cf�Ҽ=v�k����d�ď4�n5��k���}�#�C�9˹�k�Ss[x^˺tu�pvK"�q�^8zӛ����.�v��"�nM����C13� rE>�!�Z�犎��k���JH(O�Y����TT$�d����� ������Đ6��8�@�$4�4�P����l8��q$%a0!Y���l
���!8ɻH�b���$�<�BI�x�<M���LI�`^�P[6��PۦM� ���M3LRW*l{@� z����8�X��I1'��LC��d��6��6ÈM b���!��hc���u�[��� �;%d�3�/Rx�bCO�����'��x�+�b��4�[�5n���aY=d^0�s,��SN0�/��6�c�FШ.%|�2]ޜ���w���r�b���lsY���R9|g��N"œZ�I���ls̩�S|�u�o�5�oT�N�L݁׌�/ۃ��sc1�g���sZ�qX����.�Uf�gu��*.0�[�кi�ۭݸʛLD��馧�]�y���K��N����@}�	���FR�cňg7Al�ad�@l$]��Hhv��8�=NV������5�gSC .9��
8~#1 `g���-NHJw_�h���-�-
WG5�4��W�b�g �B��ƑE��ͺwXC"s$���XN����7��H��H-��[����Hj�9"bn��^ u<�����cPb�yl3"">?-���\Rp��4��2L��s���s�6:û��8�x0�o�yxE�eŔ9`kY1�3�>fX��d��l��9a�*f�Ѽ��`�		+����~���6%�b�_䫅���f��-D�}�A�c������'��h�B�2�Y<|	ɱ��7�<-$����5����1����7�!���� ���Ez�k,e�c!0NDc�&\�^�]��J�0"�Aۋ,�o����n̨�7 5 p6��T�����)�`�[�e��P{�M��RR��z}Tf9��/��<�]��#β4a�
�_  &"���w����_��̗��f᪊4�ֱ5�ML>Ŵ��= �_��C�z=���D���o�ͅ�L����7�z6(�ǁ02���fy�2�8�yH��'CF�1��D�z1`�,�C�Y+�1gg,*�ZS�� ta��o����F��(7,�\;��֮��zF�xD�kQ�$'��+����|����l8VbG�`1��z�C����BF&pj�1ߕ���W��{Jޱ�Ă����G9�ǚz���&I90�g��G1�O�
S���>5xI�|��g��K%'	:u�~H H�d��ó�x�0�2�\G^%�.�1�f�j]ۈ敛�}'��f��!�۔�f�m�7������_���I!���ڜj���~��&`����o���r�Sg��>��&0d��4�8X�J	$�����޻m: @9��V��봙ޒ��f�K��l��q�5�n1���kv���u��wFe8��C��&ng��h�N���r�;om1�������zیku��Z謦��q����P���P9X���V���tʱڽw;<n�u�D,4Tu��Ok]j6�<m�������ae��y��`9��{쏂�7��GE�:z8.����c>��l��m�r�f�4�;�>��%U尜����y뗉�t�ƵiU㴬��u��G��A7n�c���g]�n���홎E�g����a! X �$���I+$�*��J�J�+	RIa���!RY"� R#P��b�P�J��	�p9w��.���N��;�uۯ	�q�rR]1��N�덞8���0�j㮑��c�^5�9.ţ��-�{��_&���x�S��?{�����!+q�>t0����ŁD��D&�w��+���Ԙ��(q�k,Ї�ـ\��4:`b�<a+�*���@̺���/�{�3���`�Q"ǅ�D'��U&�1Xw7��1�a^(���nA��=a�}����E'�UP3<�}�!�H��V
����d6�1��8��^�&�N	b��0IϏo�5��"z!�<���}�9�E3��S�h�预U�i�;-P��>M����\j&�{Ek�"�|��O9pB*�[���X�X�݁���O�I�=aQ�N�4���x�c6b��酆o�O]y�����}�{����i��7�����˳��>��!�`�>��'Ū�Л�c��>��q� ��+/ys9��[;�Y�%4�J!��;���%�n�2��<gѐߞ���>���b��
��'�����˛�}��hQ%���^���)�f!֧�;�b#=38�W#�*��AA0te��H�4�y�hd��1"��S�����n���nt|d���R����w��;�M���ϵ��ϰ����R�A������s<
���L;���9��,3%w�Md�H�Vbb�9*kkP�Rwۮ���-o��S`�TI���\�M�CM�����k�\�L=L�p��,R�V0H�T/�gҲi��FN�{�:����˗F���*�)������
v���U��B�-�_"���
*^�W��S.���"�/��X�.�$	�ڜ��k����<����kT�Lq�J0��-_Y�9�û�u���na�zTvZ�"��\33^f��`�2��z5�e����z;�s�{�L9֛:#�����h��5N@�2���a�3J#t��S�Tm;�P�����c	��I��3Y����t�sb;�C
��o�m��0VWYX�%D#��:u<G��sE�VQ��j�����w{����+�1��;>��s34>`h�G�#�o�3e��s2���:ئk�N��Ǽ�M��m��Y�N�;�14q�t}��y��%NÜ�18��}3M�I�jo����j�:u�aN���a՜�M��S̴r'�S�>]�5�d�Ƴ�qے����r �fT3�s&v*O�
5���*��6�i�0�n4۲�i |غ�2'�A�r�i7��P1�����B7<�V��k:��%�]���&xӳ���ڿ_\h��yx�T�޾�ߵ�-���n!��Qu�#2���'��u�3_ZwLG�ܔ�A�2�L�<���LT�8��d�I:�S8���%�&Lmns9kE�*�Qb��r'��t�e��;ϝ�PV���|�B����gy7N�TS�������=�>7�����ע����hnʠ��ݶ�߮>]_yQ�**��G����խj�$����'�c-֪����/"9�\�;��\b,���?���'��L��k��@���ɦfl�u�h�XdS%�<�;v�o0<�f���5�>W������]�η�+姖�[`a6C�N�D�#����-�����0�ǚ��Y��Z>O~o���A%0�-l�:v:���f�J�t^$�Me�'������/�%�����T�rᩡ��	���D8�u�Cȱ^|I�ǎ�J��W&�3��W�ޫ�¿N�jW�t����økZ4sR�vfh�H���i:LlL�A�iP�L:�D�ED<@�8����]�����ȝt�L3m��GH�T�?i�)�>J���=�E��:|O|=�!f��,=t��1	��o���a�\����0"�V�U�6�bœ�N�m���n�h�N�#�$L9�����ΝIQ:�T����N1/o=(�ʰ�6�y��Qv�Q�����B��R�܆�;&'cZ��w�۪��Om1�u��hO��&_R�9�.�t��$pi�أ5�у3C|ȁ�W-Bq��LX(��b��I��&[�jh'�����8~�v�Rτ��}��e��b�ϼ4y۫��Y�@��o��r1cIcoI�S2ړ�D���#^J��Q7�j�fY"��Ss�Ubk�!>�31#\�U�ߴ��L.����csq|�5�T������]H�%@�,�;�1�)8O�ϻO>�~���n����*}S�m�Ů4�[!��pN��7=����n��v�GHt�q�6n@��v6�aM��;v�ým��ܵ�p��Z�Wk�d'Պ��90�k�,�\U��n-��p���a�ۢ�D�u�/p<�,�#[�.BL�.	��k��C}z��II����S�Piu8�T|��>�Cb�I�[S�ͷ�`�q�!�~3r��2�����N���$S|���Yi�5������";��;�@Tܷ9����H>����D��)�!ͫ���Ec�U�w��/���=ߝ��P@�`tp�>Z�8CI��.%0�w����9h��i�S�#L�\�w��X[hN��HK�b�D�5�%U75��t&Ȭ��S��ʏ��V���	��f���ED�3A�Q�@�=��n��}�8h6�...J�ﾋ�#��HS)0��_�����|�8,3��W�[�`qe1�=�eҘ�뉨{����~�kQ7"�>_��4�E���=��V�!�N������Qto:����N��[�n�T�;p�r� '��^mg�އ�:��>�T�W���x-+z����?m�f�h��ㇽ*[����'�Sf�oh�=�{��65����|Z��-)���0���Ƕ�`��B��}��+Kd�N�R[�I4%�Wq�u�q-}���3½�D�5��o�N��Kg�f��k^��;6�H�W�/����7&w/>$iF!��o���;@���O�����7"S�� �QDc-aRE��b���,�Qd����(�E�PPU���@F
,"0�EX���"�Da!�v�!���a���q.#Ë\��W=;�:�O�9�u��$c��0K��k#�,S!�C�5�0s�b�~�cS�̔���q1b�8�����&
��n{Λ��(9L?5��h��
(��*U�׵�-tS�]��P%\52�j�U����6e��؈�E<޲G�I��?8�Ͼ���z2_G� �����r�6)��z'��~=C�(���"f��]�S#�@l86�v�}�� ���8S&��k�nq1y�7�"3��"bz�1k�G_�'_A�1�l�!�s�[
|$Ў�)��bk(�R)�y�����O�Wz�"���:�f�*�& �ٯ� QCw_j�~6N'��5���c�i��sW]0���"�G԰Sbq7�wϗ=�ɹzn2tT�aiT�폏)w�a����b��>���<�*E43��ֽ����¦Ь@����g�&���v�>р��LE5�*lI��`z��{�̻*�[����8#�be�+�	��a1����}F9��k���9��T��2�=���%%��{ǐ1����}�_8k	�w�dxC���n�@���	f��+|�Gư�3����RS>Wh=�(`�+E�'gAP8�W�`�)��O<��.ġSxP�?7���觮�#*��=rS��9��:��F���0&n�-u�/gm��v�W:z"6�+
�Y��E��W���[\�I{�)��t�����~�����0�g��&oc`S��{߁ݷd�b8ӨlC8Si��y����>��W�d����>�8�6?�1#�#۹Z��0K	�c��1ေ��'Ɔ�Cԩ���P���OQ���.9���_P�'��)3�Ɗ����+�$�����^�dF0�7u%tFQ�j�wc|9�~=\ޔ�EP̆<`ձO�y�,�=h��l�zX�Ɇ��U���F2	�;�e�$U���{�U�\Xt�3@�n�.���n��K��������jC��:H�.j����@��#��'B��5-�C�ga3�P�ҏ*����n���W���$��G�oz5䳕bt3�̇ن_9����"���7`�U�d{q�� ��z��3�w�>9�F.��'htB"@�%-���N%��,S��H&I;��N%rL��Zғ��fR,�ʹ޽�E��~�L4��\Nz�I�}�C9ś�ǻ�_�@�çme�t�;;�ZDҹ.Y�kR��|o���*%��:V^Y��K-
��\g4\d�L��/%��u<��:`�n�z٤�J���a5�q��]�^^�Y��j��DF�R�FW(�k�}]��,�Y��t#�����ꓺb��
�$��p�P�3N������w_`���Sٔc�j�����m�D{��V[�}XO��SN*�̜������G�*�wi=2��)c+M�}��G��D&fcݮ��ƫ�c�ɜQD�V��!���F���V���f7/@��S#�L/�c_4���#Lx�dö��T�r>�cL�4�*��E,��o��/��-��4�ߟ��I��o'�*�i�V�� J��q���3���������%���4���o�k�1&)9��n�:m���y���^����ۨI���cX� �A�(nW�
W�ף�.�ݭ�<��ф�i:�l����uri�GE��;(��L<�N�\��~��ԗܸY��T��J!���@�1G���<?݄��H����Xi�����=i��e,�~����,Ҫ��S���V,�$����ȱx��a����̏��#�wI3���k�G���K������ˣh��%�'�/��I"�Q�Ae�oPb������r���V��J原Gi-�n��l�ӵ_Rǝ�׻��ޟ�c[+��@�����c���[G?��%7��^�;���뛥^��RL�?>�dA�^1v@�lD|Ϸ3���N��j����>"����!m�]MЌ��Ti�j�4y�=XK��cz�E�f�y����2t�-��W��l���ۍ�&V��>pߤ�°ep���-
���h���ϋ¼b�YO�k�j�6�I�z��E��t\�eG;�_�'���4Tx�,s	�g��$��K�cy
K��f���k-;�C��5f6\�9q[&ʝj����0Ey�x�z�v&��񺭇w���o����*�{�Fh�w}3�w��oV��?>�F���+�s+�qE�7(6
�;b��BI�'��/���{�S5�f;���>*�������"�8�c�'sټ�=9�oL�d�D�Y2g��F��qG��#�\֙!�#�!�Ei��z��1R�ڹ��j�4<����:�e^�mלy��}���"b��d���a������1D���"9���y�]�����@�Q߭�R8�K/WW8�3�JQ�4�T�U��1�e���"�V;�R�΍���(돫c��T�g������D������ոu>;&#����r��.�hD����,��ǧh�V{ȿW��&<?�{��
�����,Xv��e�::��s��}�ῒ])�5�LWyݞ:Am��c�!��s �g�Q��^�4T�I��-\���]y��2�NyC�Cݨ�<d���=�<��,{|�}�z���4	��{lo��/	sS�·��I<Ok[�I��6{,�U<��UG�������㧧^��H����3��@E�w8v�G#�f�f�a�����������}�^����N/d�nA�gi�Ӯ��P+�{Ա6p��3ƎkkO���1P��0�wg���/npE��|�Y�ݱ�ݺ�e��F��y{-���v��IK�:�����v���O&]�k&*�sۄ��8u��OJn�#m������;\f���g�b'n�xcq{qnt7\횄h5��v�.��Z;�ex.\h�n�ƣnM�=a�g��w55eC���c��8w1�="�l`6a����/cӃ�q�N|�	h�쏎��:ծ3ARb2��3�5"���R	�~��T,S�F�I��c�O��BxF9�pq�щ�8^W�����Jd.5�ƛێ�v�+&L��ȯ�4�=u�ګs����!1	�TH,�~�Hd� ""Ad�IX,
��$R(���FEQEE�+���U�5��"s���jR�ي�mt ����u��/8-�Ľ�-�b�@�ڧ�x�B*�U�>J�bb7me��Bb*
��~Y��qw��ʘ�}ݏ�F�o��+����b����(���6G�6P���$����#b�����q�������9z�<dC$���Ǳ����;v�(�!�Um&#�[8�;Y(�(�����aۻ��<5/f}Y����tݖ���N����ۼj���A3.�C8�&è�]�Fh���<�6}W�����V�����mj�}�,d9�38�r)�ٖ���,�9�;9�~|k=<����,�qʗ����g�rg�&�. �g҄����*>��N����G�m��탫��a�>q�\s��?J~�u�6�%�(�e�H��d�i�[M��9"�[��,�W'JIQDZ۱��̓pυ$x��]��=5�wR^��<0�AZ��̅kkȾ�!8��*{����.��x�#�yՔ�*,U��^���G�dڱ��"�~C>jN������l��%�D�j��Sk�xN�%�*-V���Ih���¨���Fe��t{EE%�̓ѣ��Dk�b��͞o����N��`�9�:4��ޗ���FU�>��3�q�֝��_9�,���"�H�I_My��̱��q���y��D����ZPG/^�v��Ii>�����׼<�izM�c�7'+c}?_��~v���D�I+�aW.�x��"��Y�R�1�=���hV�epۦ�ߗ,©�8�!�(:F���L�s��U�q���|�y���[8�P��zDI8ƴ@��r�9H��&t�9�����5��mD-�N�AQ~+}�&�k%{Um�k�JP��d�'��76�ޟ�5`�v�n ���b�k�ڴK�9F-��ܱ��O=�;y�ێl�Sp�N�T���1�m��Ve7�+�L��){7Y(��,��xҝj6���s��%]7ۇ�k�ÿ�K3`�6�*vvGmԫ�5@��:�Ci����5y�Y�M���Q��yl��}<?��xj���c�滾L�Xٟ8��QvY{%�n7��-����O���Ke���ޮxװ��@��r���6#̰���x���W�ѩ���UV�hW�v�Q�N�)�J�6Y�T��=NH�E�<I4��4��7�Z��W��=�7sz�^�D����ת����y���%���/�Ϸ�Β�!�:٪w��T�Յƽ�7�?k��Q�b�V����W����a^}�����md�d�����՞ߧ<�m�	�dy�O�6񫙞1;�a|^��Ac���a��Q�O�|Zhz�i�ߝ��Ǽy��]�a5=�N]��i�y;�q�G��^d����5^6��|oyа����e�{����yc��1�(R�FF�EF�δ��U�J,�H��1�c�Y�]i:r��YϣOC��K����e_/)�9��f�G�,�1D�h��c�����y�+!l�޽}6g~�>ُ����p� 3�c�A�nֺL�z��b}Fg4�S�W���o�w�巰�,xI��i�q<$8N�+�bګ*�7�"��Ʃ�]۽QN�̔#�k=�S�}k�B�.'x���vu�v��eM�8z68��7�Y�|���y6��8������ņҜL����.�'����j#���,?k��O��p�Z���a}Ïn��h�*#��A�X��	���P`-��f�R���������� ��  s�\Ů�nxN9I��	E, ,�ZW-W�W��8��Vkz�d���Z�%�V����W'�Ź�qD���yL��q9�Fs�䢸���I�������������s��L��z��8�h�Z�K���k<o}Y/�#j�1�\%����8�[Y�[���>�|�7V0�v3$�d�up��>�zS��X�7Lk�T���/+n����N��,|��MFa=)$��
(��������wNM2fT�t���t�4xStL1|7o�ظk������w��W��l*�94�E/t��9��v0�i�Y1���k���b������m���u��0�����ho��=��Vx����9��w��$�.��\y��a�\�/:3��Y}{^�|�%K~��Z&��?g� ��S����e�nPU���k�x�ۻP��<�����n�cYϿ(	���:���L;��ۼ���h�:�.�oe�9z����n�g�*I؈z����'<*Ǟ��w��?2�,kط�!���s}�Os��SRɦ���F���^J߶u�f;��<���������O�o{֩a��͟[��{�A���;u q�Q�q���.3���ы�)���}��7կ�H����R*�X(��RH(
��P�E� ��%���o�F|�;:����/0�����Rm��f��;�&�|�z���|h�ث�c�/��4�V5<4<@���*�
��	�ד~��.M�Z��I*�܏$���w��A"-��ϴTj���3�
}Ky�~��7+]�K/3�;d�r�;����ק�d��	�cmpc�x�8��r���6���wH��߇=�Vش���;0���}5�\�yI*+��hqH%rV��Ǫ�g��院H�cא̓]G	�c�~��ȏM����φ�1c�Q�n�)^���,��$�!{"j�i��3C��VDw�}���M4&H����"��J���b�mY.�:���Ƥzo-��#1گ��V���\;DѪ��j���tUE ��ʝ��ՠ���yH��[q��t:A6rk���n�tTV��=�l��^š��؊ �F�V;0t���U��w���H��.�q�+�w�%�5���+6�xa����'�t7å��.�Ȧ}���3�D�C�	4������d�ه�l���j�������;�5l��������^4kJk�rn��7��AIc@�D�c@���e��LF���3��:����t�~��U�g��x����c��'����ܻ>�A������%��p�:i<u�&I�i���.XTX�Y%�{!��O��̫2���,�XYq��:�'_viϬţ"(p��*೵7���"p#��Bq��-����<�Y��O�L�Y[��1�=���i��f��ʡ�3��i��62v�K��1}Wcd���2�	�.-���wK�����[w�d�ɶ�<v��$��ޛ��3g��}�����R�:D�Qӻh�,�.z�ٜb���D�F�hP'v"PȄ'I$��a�n�m�¯aaY��u�7��N�Q��g��ʬєY�'^��M����,T�LQ_%��|�Ez�]�m����eg���f�z����7-�U3f4�*EXΕ�\�>�v�ʴ�\��@�H����±��W�����������l��,3:����h���*4������E_O;��r؛���>.慻-��}*&ɾѝ1��zm�k�:�O�lYj�mԤ��7U���J~a��ie�ʫ�d��M�.�h�h�×��YEMu���˖购�|yv�M"��mkeTc݌���N�/=���ւ�Nun��W>@����.�z�]��G2<v�\��c�h��]�z�t�bT@��[����M^{�뙬�&t��n�$���=��Z҉����oO&CцW��3w��h�1t`�����cNj+vIOG���m��k��tY��g�dkJ��4�xRt<Y�B͟"*s��\������m�9�[�i�o�:';"�k�&�yu�꘻�ݱ�[n���6���0�'�:72����3i%f&�h�F�g�������]x�N�zɞ��^���Ɔ�B&*�K�)���J:�0�y\�3��ι,S
�kl�T$AG*v�/{��B,(�mx��;��^��^劔���y��c}xA��؋.��H��69�����#v��A�����{�z���|���φf.��:�%5#�T���;�_]:��ѷ�T�d����#�w$M3��Mtͱ&���N��zW�r�!����|� �qb����[B�Aȣ���bم�,�^�-�)^^��L:�}��u���(���Er�1u<��(�hn�d�����Q��I2�5�/�.�9eUO�&�]n�I���I���`�A��>5�sm��Y0��j<�ՎΏ
�a�N��˓G'(c���xz�\��c���R�G+�9�G��|i�]F�d������=��t�i$�.�#�o�̖�k&5�U'u�Ǣ�'n�n��Û�F��ǝ:�;s}+V^�;�s�6T3���{��jvXIͣa�?Q��AC���/�G��������ŉ�����r�o����>�BM �=~hǛ�]�z��~^�=�lz��#R��}�G���=�����ᨄ�����Ii_,{��y<s�9��7wi�V��Jwdѻ�aX����
�����4x2Y�˽�%g?n/N;r���T�ɬ����4t�5L}���*ȴ�W�z{p��7snQ��N�__�����������3�7����h�=
��V�sz�ȼ{�kw�zұ��yû����;��s�g8j��7�(��U��z:��/���b�9���9�qq[��۩��n��ۼOc�����wl����3\��M��xn��[�4p�������lu���؍E���q�s=��n[��m�o+�x�!��,�c;�qƻ��p:��9[\ڞ�۝�j=�`��WtU����ڵ�GM7�Nݞ��sY��r��6��ձ�����uOh�<u�F�����E[9��k/Q{j�cqc�:�9؍��I868ׇcp���2�ݎ�k�:w+ls�/�#����<\v;g{Ov��V��-��[�N�3���q]un�=��t��c��]�>H)(,!
�*
�I��Ea"���w������M#<�ע�ɉ�8��@��� �m�&1؝n�pv��<���E�oo.��7�p$����m�����1x~ ~{����x �D�).�{&~���N�l�-�qM��ͫ4����%�֔��q�7�k.#�{����i�w"��?���;��:Z<������1�v�1z���fƙ� ��j(v���D�IS#��l��1�/,�	�˼o^;?ciS�.�r�l�x�[��h�N��c����/S�C���m��C�˗xR4UGS��V�[��>���L�ba�����	ӌa���RYD���8�\�vz0����Gho��K3��Ǉ�,��@���e��%���2�o���fϣA�˶���Ừ�F+J��xß;p�X�$Uic]4�^��~�y4~��`d"��ܿTO�+|w�d�a{�J���I"���s>ɥ�Q���K�z*��m#������o��\��`�)���A��3%���YT5��޺F���k��65��V���O�uh���T_�̽ގ2*D���FE��#u�;p���[�XgfM5�"������+�SG��g�����SU��%0g��El�;�����	�O~� E�{�EF�z|���I���TP+��#vR�E����&u�-�;M��C��\��:H�՚�[�_=&��cq�

͸��IQ|5%M>g�
�v��/�K�����UI�}������6�y���,�Zm�g�ᥦ|�N�ǌ��x�g�ʙUf�6ؚ�L�� �L���2l��XB|S�^3����۶+u�;U��=�ٹ������8�#���6+<vj^4����߿�����]d���E1$:NI�l�/�YP*��b�VI֠�3Q��U	�G���>��\���sSQ�ux�v��'M��+j�Rt�B�#�n���g�����8�NZeE�{��'0л�3|���i$�B t�4��I�BIYIRu��"$�m-��{���fK�Wx5���]��ۯo�	���v�-���s.����E��c�Q�~���k��d���H���xײܩe��B�wU��s#x��(�)���z��.T��H߶�M��[�s(��یW}���,���Q���¶�L�����jn�����VVM�_�_�P�}y���g*�ьy'Tm����L6�֓%�=kg���߽#s6��h��ᮌ̲v�*�Ml�Ga3�r���fz5�[$`�۾�KX�3S��I��&g����be�D[{{��_rڿ���A ����Vؚ_���3��U[y�Lf��o�����.���6���
�i�^�I9�g���.�{ɣ�7R.����v�wᣆ�|��2���3a��,ڦrjj�8x��U5�3�$����0\�����8��}��y��y]�B�\��(�V3$�O	:(P�p�l6Amҝ{:�gܝ-=\�/���pYa�-CG��#��N�a�����}6z�Y&a$3}$ϒJ2ǅ����9Q�M�a�oⲣ�-��������F�BFdic.9���y�Gzi�VW�%�[5�V&�i���K�9M�r�qJ��R��Iw\���w/�#�!i�]��%�c�#�4m����.�,�q��j���ٹS�l��+֛DS��q�w�w����e�*.��-�fu�e$�|Z~gs���nK�/zp�i��\S�Y�&������?�H��7z�$�n��4ua��5���e�]5�w�ʉ9��?���;ѓ���O�;\-f�Kh�U˻���x�F�k�"��
|�2o;aDF���/����M�����W�|�!�l��V�>�÷u�b����|�$a[|�/!���d�CU����D���Ϲ��C�@��}�e�H˼d����h�L�_�mO?���{��c��x����2K�ʜv�')U�[j����f��-u_t_DX��3<�I*��5�2��o����ש��q��/�I΅��|��3�k�-抟�_/үc
QY�j�}|������/`v-Z�o�]d�#����>�p��y�r`{-�2WJ��S���z$.NÆ�׻T�RͰ��=�/Eq�9۞���^�W=}A�N�G��'���읝�����1�J�+s�����~��_<+[ȝ������|�����7O��H�U؟��eד{��-Ƨ�T�M��x���ͦ�O��{���O��xe���m�c����s���w�����)"��T��"�a)K`��"�z{�t;�y��gQG���!�4���.��7�2g=��iX5=�����34�R��;���+��X�&�ns��kjh�R2�ZUkJY%�\�*����OLw�8��E7{u����槃�.4
J��ҫ��0��wK���w���+p�i݅I0���b=�W�+jgͫ����l>����=�f{7��w�}�|����9Ǧ<_�:\z�N�֘���E_=|�~������Qޗ��DNt��+�?��[Fq�H�&+q�����UFc�+|q�*���T:LYBVg��I�����aw��r���G�T��^�d��3g��q����q� ���c�+�l�����$&��|�0<�y�Ahv�{�.x����##`Ơ�urh{�om�,U��\񞵸���s{u�l<V��k�.܍e�7M5��竇r]a��'�Xp�Ū�;]�~���x|ቔ餹��*5��,͌��6=�[αEc{�Rt]�,�a^���$�#�����'��c�,�}3vP�S���=�K�=o��S��n�i��ֳp���7}�UB@��--�O�VW�~��,ť������й���wu������'2���l�c�_kvV�D�J���㤶���/L��+Z��bI.%����>4�߲�0T8�:;��7_9��;xO�{�'��4��f�y3�/��A�<c`��Ϩy�����
�H�H"�R�-^�}�m㼴ô�GSo����Ru��:�Nv�x�lNn�DWL�C��'t�0�_x������\��y.�|�9�gɵ��lUZ�Cdǹ�^$L}껖�m�{2Z��2�F�1��=��O���4��n�%V9��κ�<�/\���]4ɡ�����m���%]OK�sJ�,�eJf�򓘞�L��;M.`��j2w)T��{�w�����YX�&7��rL*
�Lf��|����;��b��Ï2�2y㪖=?O�/	]aj�����N��z{�&���_s�i:�en�#�~c[��̳��WE"�	l��<f���.]C�т�f&d�i����70�%�p�]����T��81�*��QA<��c;�.5�0�Y�L݌ƻ�~�;��P������l�D��@�Nc��K���y%�y�35`�q��Cz�,�x�(�#爢�k'�&3����rv�i�s�i�Ό�:$}�D:��{g�/P�b����յ�N��W�]	�5�z3�]igu���� �+ͅ5�k3D���L��7����k�m��J�nxzy���vI�>����^��,dM�ey��õ��\ǶV?��=}��ܟ�,U��i����O�m��e|�BwP)PFFQ�H6��K<QJ��{��k��M^rӖ[Ǯ�8�j��Ș���<�*b�]�s"[wM�<;�b9QyR6[8�{�����8M��PT�o*Z��*���<-L,9s�G=�B�I�"�<-�gw7h�&��7ٜi���߫vuX�ZY��J~��9��m�6��u�I^����d���7N����L7鏙\�w����b�����ƾ�쬋#ʦJ��Ɠi�U�l1��?�캿;�����
�t)��$���<�$�X�[�4zoʘ��ˎ���]�����ϛ�aeu��"	S;��/M�;��QtD��~0Z۩Ң��wJ��H�����x���\bgHi$��k���t�I�o'u�OD��)�S�n��ߞ#SB����6i2i����{S����{H�����r��Id�p#ul7�� ~��v��jI�xN��:�0��*�u��]]�k�!yw$���sx��,��ݭG�����S�)E�����|C��DﳔGa��Tf���d�̼�cP�47�qA�דz�8c�7$�hn(H�꾙&�����>�����m-���y�w��72.!�-�8δ�VsTf�T�p�y,G7��4ӝt��e^$�Ou� �ɤ$��nW=s{����y�v��Q��=|ͮ��]��96����o��k{�8sx�q`�-���>�l
sÞ6|�����e�c�A���ݚ�s��zm����{�§�<�l�v��v:^8�~��3��),H8��f���o����d�N�����S����p̪"�ɕ���|���cٱN�넧P��#�8��x�s�Ի�6��x��=�-q�bz�փ�����p�.�4���2vn��<��5	�6ڍm�Id��|v��Y۠��v�v�9`����Fzy�ۤCWA⹭�&���eݪNva���g&;r����[��{V�������l����J��U�ݻs;h9m�b���8�e�[tp�K����Ob��ˤ5�±	F3Cn�	��l�ۢ$�5���ۛf�Övͻ�;��z4V-�k�j��7r���H;�N��=@�Bb|��pՂ�G!=i�6f�E�W4�q��*@U��dV"Ȳ,FE�
�0Pk9��.���(��C*�H�����;v뮋��qt�w;u��6�/������Of��
�k.�t�g)-�n�(�A�b���R�j�=��L�Kd�-��X<���t�����=�/	�#�1k�4���<61�1#�-�첋B�^c����]���d�3a�z��<d�����#\��o}Ԟ�V�ݸ�$�`WU�v7�0�wXn�p�j/�{	ű�m���d�w��I�l�g�fˉ�K�ӳ]�t�f	DtI:-��vk<z�}�Q��F�&�wu��筝�u9�2����-<w5[�6��t:�����f@�0ś�G{�K;�,I�ã����C"21�D� �	21j�ko��yvG����Y�n��	&�Ҷ۔:�=P_���;?�=O\�`y�ɢ��ˤCH�Xʢ�*���3�+�x�P;�l�v&IFP�A��H��94<���v�j!�ѻ)�!���yP���[����#Ï�-��IH�v��1�����q���oV���N�]{���<g}��/��Q]��I����ꪣb�$�Y�x�g��=1M��kEJ�]�]Y�������^��xE?a�E18�6`�`��yU:�w�$[�:��H��S��c=��ط�F�6u�9m��渧|��tE"8�8�R�x��`n��*ɖ�n���cϾU��Տ_7��[�9�<�K�T�w���0�����m�l6�ig������K{�]o;�Gma��-�`�y�rn5�zfV��B��k��na�z:βvg�/���JQ�$����!�i��h�����z�ڋ��3�lIw6�[k�架�޷�r����C�I��%�ܘ�����Fⵎ���3]���oӂdj�{�a$��I��汕�ǿ(b�(��N�6��#6�i��'RUv�DC��?�,��^v.�|Vq���^�3�N��ck�w��{:�0�og�ω�~4��`�4uݥ˾�,�D��:W����r5`"QRY!U�/y>�mNcYQv"������ړ��%�ٝ:����=%;�yw�孼Kޗ����[#�'xIu~2���N{Ν9Ŝo��y��KQF룏Lm��Q]���Q'��p�fcY�[Fmv^�'u:va��IE�\[����������TRVԪ��DBx(�",]�z�&�k��Z)�����X�����5=�ۘ)�|2\t�TP�6�~�<�7�O����ɕ�l�cCu"DM����&K=��S}¬9���&�p��i����8�T>߲F�Fwʉly�ڶխz����z�	贳&%E������~H��(6�L]��ä��e
*��E��7*;͹�����̪�/��W&^�Z&4�C�<xN�����뫘<���o[��ӛ�|�}�p�rթ�X�{�=mRn3i~2�ltz�q�����¹�w�,{�`��D*"����	�F�V�:�a5���1�n�fQ��Sg�G�Ϊ)t�rD�Q���:Nc0��ag��^����d�3%�nz:E��{FcZ$x���[�5��C�:z;�ͧ�}��";9JN�b��Q�C�����(�I}����|�e�=�ϳ��y|�Gr�ušWgk�m��X�z.\Z܌<�{7Tp����mecR�q+����]�;	�E��+p���c�O�XO7N��"�3͗X�&���|�{$�p��jٱ����Gug��LA�ǆ$�M�m���øӟn^�}��_����b��<{-߉�󳯑U����T��P���=�k��ir�Kٳ���Q���B�I���.��b�.�y���sj{�i$��zn�4fWX�zk��d�D	��Ne��^����PѤ�S�G�g:JrN[xc$��q��v,�Ev.N�c���[e[�V{��"'%ڙ;`�D�{1�,aj�ao;��^�����,�F�іv���'�μ.�zA뻹=��;[�C�K���a�dz(�a����ʘ�O	������:��g׳[�EYKGg�o~x�}�|f{F2z�2�F?��;��?4N���g�K����W��֓D��,�݄ �o>���{���1q�]-�#{�.��;��4zJĐ�v��<Ԝ~�_�O�&�qz���3��C�DI^���<#��RƩ
S������n��Z����=>��$1e�Yq).��/���\0�5���ߒ�˶��8���23�-�)���I+���U��G��a[�9����u����A��(
�
H�� (��|�4_���l��_yۉ#*��&4�6�K�+��Me�K�Li�,���C}nv�o�t��;;@��t�<BN��s�*��8ϴ�fɢ+'�|�(�Ϸ���&Ǎ좈�쮝(��0��{�x#4o�����	x����#�m6�;��Bgw�7OX����ǟ�m����	�L�78z�	p�l��4�o��8������7=��˄o6x�:R
d�W�}㾌j&y�Yu�2='���ޏ3$�G�����tY�E[��}��_u�(��e�"M�4���j�$�����=��>���*[�Y]����<��O,9�b{��Ќ�0Y�y����y�g���֓c=V�A���댬a�,O5�%ձmXlnN�:ŷ\��ѕ�l�;r�nx��6�:r(&��u�*֢m���D#���Gĥm�N��U������e�e{,�v�������_����8�+����ڙ$q��1�v�k~���ys��J�=�1����4�DǬ�CUN���I9�ōj�]��9�����Y#�
9EԿH���-F)����p��˝֑懴�	�'�fv���y��}M�X�X�t��u�T�"S�ӌ�E�����Ec�Jd���{<��ӣ��>��$�#���1l't��/\��Q���6�W���ԏzO:y;�z��J;p�8h�����]�Fz�����T\}�3
H2yL�Ww���"`U,ξ�k�����H��%�g��J�y�R;����Y��e�*<��Y����q3�v�&3��2�OJ��+kS$�XR�-"���E�0�i$�Ct�{�h���5ñY�acj�(}�����D3���ަ6*W!d���k�[�9��wјx�i��g�����j�0�9���ܩ�&�Lzk*$���CA��ZZS��w�Z2+��D����ob�ƞ�y��Ke3Jͫ��!lqħ�S��EVxK	뻆~:��j����З��$GІ@B�@-���+�z=��z5w�w1�_s��L���h�۾�4�����IǑ���jt���d���&OS�
G�ފ�|I�Ƙ�����fd6�k�j�79�����a����
.�!�|��h���Lm�oك^��8�[�5���kz�"n6!K�BK+�nfӂ��v]"틒��ݰy�'iK��l��b���;-���\��h����!��6 �:@��D,��O^�<�<�9�{���σ���o��,.�Y�%7�/N.&��{�[�l���S:���]b}�_DO�*尧i-�g�d��=�{G��X��P�՞���R�Տ
�����=��t�_Ϫ��oy�_���5V��p�"�0;D���Ōb-��g����V���L&9���e���׆�K�|^<S�#Pݟ����cq�MtY�(8]T�����W���=|zs��4���j�y����q�+p���ayQʦƗ�U~vI\7���&k�����I?;��}�oL��"�
(���	��C˫]�wϳ+4���)�Z�y�I?��cZ��}��e���O�m$��/3�i�+2�WK������es�P�K�Ot=������_*NMR��o��<�{#�3�Fs�]	�[|�(޲8R��#Q����;�ݕ��z,i���*ݪ
V
�B�h��ard���ˁ��d67\���i�q��^��y��c��,}��_���t�gkf�|��n��H��'*�:�+Hs��-��X���^jxަ��z!��a�)��"�Zѕ��y+:�Jnoa�H�nI���x�(��n��������6�r����{����)h<=K2����j/�u�u[*8�lϖz˯N^,��q.�:q��a뫢k�u9TUo��x�}i����w*�'�3%���"�]�̲��{]��� �?zVJG7�
J_!��m�ꙙ	�Y=��R�5vQ�4^;W�,�z�1�>�.�j��y�ϸH�{���oPi�ݞ�A^���o�p}�C���<��r��a

�!�L��y��,f��h��7���3n{�XW���¦�����x�>��C|n/uY��7�qg�'�J�z�����ln�.ˣӳ�`���o��)���:��,��"O��2��j�3�����s����"�W{"�EӞ�۫��Z�~	��㭪������	m��.W�=�8mq`Cf����Q��l6և1�ȖٱY9���F���<q8y"G^yÔ��[�[+�#o("��Ν�A��x�qy��[u�	:3ϯۇ�[�������v{x�y;i���>/nar�>�3��g��q�`�5�7o:K��!\��z���+�
�0�]��m6�`�iP�;���\��r�m���J���܆��q�]��:ݧ�a����'ےݼ�	���δV�᳇3�s�*n�:�y��P䥺L]<�6!���.����|�)��B�c�����P�)�}�p��y[�Wї�nę�㧕�F���m�ϭl������{��c����V���SeUN���zw%u��Usk�<WC��;�<W�~��#���1Lfz�"���������O��{�Ԟ�t�Ϩګ'ڨ��灊X�$j��0좶��=�eݎ�H������j��ۼv�ߋG���,�<;8�:��%�'��Fߞ<=��u���۽���Ԛ\i1�ke��VF|��X��=�RϓO�-������{I:���?6�o˯����C���HϷ��:�3L���������#/���Z���.��%�Ukoŗi�X*+�m�:B�ҵ��h����.a48AI�G��߻H�X�/Q>�:������x�/Y�ڳ�T�I�s�!�c��1�R�~������I���"=��x��o;qB�k���;l!f�Ie!���?��CP�UcU�a�t:�$An�[�����	)dS�l-�8�ػ�0���ʧ��=�y�v��I�*��cϏ��q�oN���Jfӽ
(�+����U�):H�{��q��u�,�ô{������5k�:r�d����m�V��y2v�Iӕ�Ŋw���F>��XY�=������֟BB�+D�$�*�a���|��~Tı�Gu�,��N�W<p��;騻�T0����Q�[��#Uv��f����W����av�H�r=Z.��c-Cv/$�����k+J$���M��y�T�X����0b��-c���i`AA"Zb��u�s5���Co3�0�F��0��xę�Pt�N9v�L��8��=X0����.[�:��;3���+Tw���ҍ���Y�VV�M�`��s>�;m��+�4�����{[�r{m��)D煉%ǭ�vn�Ղ�<Ƿ�S�h0�o�fçNL�=7Bj��o���^α��z��'x���I,�����Ŭc]f^���I�2�jc�T�-l���P��1\�S���7���ƞ��L�\OF;��wy4Y�q�0�4e�a���q�=��#��n�5�����[�t.�N�����F��t�a�0k�Q[my�jX7�P��D43�>��"8����in�q�EW=G��#nƗ�t�Ȭdk�s�����#�Sg7��ڒK|;�3ޞC�סڟ��?<��y��^���Cf����~��n��WVwO���uǴ�i�M�ש;�=��3�.=;��������z�N߳��O�$W9���v��wu��dF@����ӘaW�f���V��ީ~T���}��Nֆ���ѓg�����ٺy��47U�Y�S�;��pQ�͆�� ��f�z-����%�oU��n�Jj.�7u�^�^;���0�w�%��M$�E��/7�2N�%��c���AN-.��[�F��/p���d�˛3��ݫ�}B'�:��ߌ3xa�g��W_J*�t�zrY�b�D��K�r�惺�F"Yw�gcQ"Me��$�Tl�̼��蚊rHCe��so2���m
`� P�P�.	�8�v�!��7mgv;l`M;2+����Gc�m�\[c���n:qNkv���]��%�vw-�G�2����1Q��/6����s���-P���K�H�Df����P_�U8���oxo6`�.������7�y�k��P#��X�'V6ߛ~j��Q�j�1ɕ�⳩�r>�Q�]t����쓤'Z�$��ѿu��JU�cee�u�Y1^�uLZ��I,z�r�-��h�������y=�o�M�U67zْ1�ܧ�슊�2ǭ�:�cOjԝQ����#��ٙtmi���I9'U��>�n�l'8�4�Y�t�Z���[
�0�Z[5�[h���uqvg�W7���{�a�W���]V|��іDwp�hf8�kw�hK*�m�TO���t!���5�#	�ajjA�ϯ�����zx`X�~yz9=��ޱ��;� �Z�&d&yg��9���d��o�vԸE7��jB����ۛ��y;s�Lr��
�4�3�����=ι�����q�`�-�I��Z��3NBO^��<8��ە��[���{�+/���4�ʬ��+V��R�'�u�8�3����{��I�ښ���}x�<0������G�¬���{ޞ�ޛ����>H�#������:�:Ne�ޛ~�#�����x9Q�kH�,��ܓ�?6��c	����"u���l��6[�E{������Q��3����Ӥr�,��楐��H��c�PFQ�{̒cg��<�p�lQ4{~���_�tꋸFp�]
�V�c��o����=/���&2f��7�?�\�SF�H����4�k7��C���~�w��C��J���Cxz��oYd�?��&��S��c�[O�[��aYF^b�y��/��1)�֑�8�Om�x��ojJ��\�3�m�}�>⋶�z����������5��K��}Gh����vq��K/l�L���Y�w����f$ xI-3����ٙ�!�¸ki+eų��ӧ�p��q�ίc���S����<<�'S���#	,�ustMΡ;�.f6i�RK����6/�L�8�E�p=욵�k���w����9~w�+̣�Yc�?�e��	ӧ�VK��VY�t=H��ԇ�ڇ�M����vV��q�앥�"џ^{�&C�fb$V���I[���{]�	ŭ�O1��{���L�j�5����٫�M��j�������R=���4u�S؝&*t�\_|�4e�3+�%�s>�EK}�7I��fi�7{�d�ُ�IP*:��t�]���]���w��W�H�P&6ۃ4<!3�'u�6�*��sz��7�cOg$��/Z�7r\F�bD��~�Ol�Y�d��gԯ�r�g&��͘v��O�r�q���U�I~<o}��$��]�{-���ۙ�'ټ�-�ލfK�m�VL�gH�-.��^F5��������J����>%q-�����\kY8��|�Y!�uYP���=�*i�lԺ��bdhdOU�N�N�����>����mQ1���B���x�u_�OC����4>Ó�/L�V�t����;dd.0���4;`�au�KF�T'2&F�9��|���d�JZ+F+i*r��d�g�����U��J&%���T������
��^��7*��QpNf�I����v+�}�6�⤯l�u1�=?x�}�5�C��x��=֥���������;�?���7�����J̅����cB{��������u��e�����;�&ȉA 㭉��`݃v��*���\x7*ݍ�fĎ��n�gE�S:!'Ol��4��������8�$�ۇfŶ��Vk�:N�I�wL�{p���A[�t?���i��Ѯl���Xz#�QՊ�:����u1w����<��P�sb}%S���:�6���ߛ�b���G���쨮yxxfB��U�$Tpe�F�լ�����5U��&"��f߯�<z#|�%4��ʚ]7��/f��o[��&	���mL^+wu���hܯ=���h�{��PԹ,d����Xn���h���L��Y���w���^��՝��<4�d��Z�R�?��|sϢ6�M��͉ʘM�ra�z܈��m�Zwy(s�8��V*��Ѥ���6k��]�}�oFG��WI�kP�l��*�9N5,�kPӮdN��ٌ�oG�kӏ)B�Y��ʿ3�
4KDR�jn��ީ2Ls��=ݿ�����h�r��Ǡht�3�P�"q���vx�2ۯw��+��X�y\�u@��;�$����әα�;�)QRI�Ǔi�s��V�/U��,��
��*~�Ϲ������5#Sմ]��~����,��gK�0Nz���� �׹�g�d��:�T��ꕫB�����춒�g��1�5zD���&5�T��Z�1Fd�W�f_EBIi)�d�ɯ7L�#J'U�GD�f���nl�Q�t�oo�4ݜ���Q�+�����ty����o�����|?�~�TQ��
���Q
(���񾓼.�� �|^�Q�~f��&TDEI�"H��ڳ��7R@1�!=�a$$H�"B0����U\�bT,&(��Bz2 E�BI!�J$_� ��UT.�B)��EL (�DlA �#D$��)�RM3$?S6�>�����ORt�C�p����DE�@T5Jʪn��ݖ�,th�@僽�G�<(޺o���L����c�������������g���Q��.���3��hѶu����ٝ�O��lM���g���.�3����Q�`tl��c?$~�>k����$`���P�IO����.:|���0[��ZB�>aWm9�_���.�
ǗѰ�W��W�t�3����� �!��_d�C����C�d{aCg��1�E-OY$1�4���!��V�0�[�V;��\���Nv8Z��
;1��	qD�UB�F�T�"(�R
	 `� )`� `) ��$X
DH"1	@�RXI	�H,���(AL� R(0C��Q�� T`# Tb�q.��	L��i���w�0	�i�4��(
!yE��!-��&�@a�5��r�q����m�vi�W��]�N���*������R����u�Q,�h�iՇ(\����V��hl.��1W���s����y�0=Ɛ��s�w]Ŷ;��h�21�t�*�o5�! ��v��T���Z��.�#F�3G�gvA��xrZ� !� �!��}rRsO)��l�����B��H�.�΅AD/o
�F<�hJ�\���D  P��4�L���0C ,C6�Jh�~'U�����95���j``g!q'��~�����%�FGW'~`�~"p U��0G��w�����f�.}=L���#��,��mT�w��$��x1^%'i�xs��h@Q	ϣ��!iHC���v�� �!Oyv<K�=��.}����a�7.���/oa)Turuo�KMA��+m��Z��OIі��+��\�cE�oԗ<�x��=0��Q]��QhC�.�jg��QA��۷I�'@��C9HVy*Pj:���jSH�(�Պuv[C�dR<t``�t���pirU������~��I�88�s$˗���R>�+����p��]��BB.���