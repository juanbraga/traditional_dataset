BZh91AY&SY�A	� �߀Px���g߰����P>]����q-�B�ۄ�)��D��OI�zj z�h��Bi�� h      �E=I� h�     hɉ�	���0 �`�0�H�4�������⧵� ���25=6���R��,��\�+=���"Y����H�g~�� 9�������*�B.d!�0괃��,ZL*��Yᑫ��ޤ� �1Yn�c�������8����" 8"����E�(�a�Zc�r5B��l��d���뚷�%/HC7׶��_��4�B�-V�\�[��56���V��g,Z˜@��$��K�$9�u��}<nUi�ϑČ8c���H���t"�yk��i<�i.�K&ȲZ`>ZC3�:�3^�m�ȗF�2r�^�,e�� :���aLh���LeB��t&�Di�H��i�������{l����"Z��,kBr&�{c��A���$� )E8������m|!�..���5r���r�Q� �D��	�eP�p"x��㕰�c�zh��=ڧL@���P�Kc�~SG�4�(�f>K��d�|�b�m�X3��&U�B<��>�R!M$�wۜ���S-��4H�#�ȳ�u(nѼ:@9�(���R�A�o��mz:���Ն���N���CoR��J%�	�����]&a��!�|�|5d�2L4�d˷���<'�
hHb�L�R���e�I��R0Ex&��R��h��D�
0���c���֫s��.&'>&��4�tf��Ime��0�]��Q�8.�t��$5��h`󐉘�Ѹa߇�q���}�L�}��=t�����V��h1E:*��4?u�է9:����Kж�Ij�
�a����w�Cs�#ŗV�R`�X��RB<�b�$ȷ�����\VGi�̚b��+aQZ�ImQ���VO�����^�����5�w��0��\%C�fOIuD��!���ْ���.�}�'F(z�v�ZJ�wv���<=Z��gv�Te��6�p���40d��G�=�.ǒEh�z�xx��Ӡ�'�
C|�$f1$�6�� �P]s�R2Ϧ]@�i"ׄ��)|Ժ!�ĒA@��� FK����B�h�7��.�x���Sz�(��#L��}ЦAe0 �r�E�h���I�D��.9���ݲ��c��
�ӭ3���H�
(!4�