BZh91AY&SYy�� ߀Py����߰����`p�s��%K��E�F�d56�x��di�  4S�$
���������h 2i�# `F&��4� �S"�J~��觔 ڃ�4 �  z��dɦ�L����0Fh� ��S�)�&�Oԁ�<�����hѦM6�� 3�@m
� �Q�}� 4V$��¯���"x��3�{k>ꈎD\�!:`&�8����y}�-`6��B��	���M &FKp1H��X���Ǌ�S�K۞���(�m��m�.N
�J�a(���̉#$�F
i�)N�2�T� r��ٻ%��L���F��hOzq�,�dh�IF68)ۼA�%iTD�ʂ�fv���E?,�����=��@$���4x�7�VO?g��e		u�SX`�Ou��Bu���S:ifv�.�(9�J{r200"���;���w�
ì!c��;6�x���$F;=ý̴˖d�Hh]h#wXI������8�"w������ݦ��kL5VӚ�@�Z��fW�Q�TC[^K�UNA���#G5�YPƃ���Ƿ��>��>H
���~l��;��2Pva}�!��8�e9�v���C�����Su.�	(��A�y����];Փ��I4���>��Uk�9̩ך�uZ�_+&i�Q�@r��&6��g�g�ȑӅr�I�,�.A���v2�����
�z�ZWwEF�����܊���V[)ش�6h��lH>��F�@l��_��8޳MZO|�!�fO�61����n��[�Z��y�o�v�!ƒ\�HH1����'��]X�E_Z&����x-7��Z1�1$�0�(H�������b"�0B�`T��Cd�?�gR�&�7ac�4�EMT̎�l=4K��X��X����>�P��M�O�]A=�?*�]}�ݍ/ݗ�9vo�g���s?�>o��[=�������8;�!ף��i��Y��%�S�!�\�Nߔ�Q\[ȕ!&��$~1���t
�~5	��Z,M��a4/�!Q��]����N��W`*cܝ��g˞��gj��(S^(��*H����hǮ|�hT̡U�-�jU�X�>,Qd�g����#�*A2#0/!��B|�EYb�Ɔuġn�0�I��ĩ�	@H
E3$����B\�2��1��t-Y�'�OK	��I��9�/�������P�*Y��P"b��ZP����80cZg!���J���(ϧaLq|U����zCn�Dr,��dի�$UkLvP��|x��4�R�郔�2r��:J��(*uTr��Z6�#��Pb-�< �n����b�1A	$l(�������mߧ���Ie�憌HA�)/E��t؉�z�+@��٤c���JXc��}�z��Z��$tr��sn�LX*�>��2o�;���;�4и"�Qd ﷳ��W4���r�[&0I��p2.	`q���hD����z\���nՖ�9<��80� ӱ�Xfg�ô�F�
ƣ���N@��a�@���d��Z�lۼ�ـܡcFq`T���IN&8����	
�Y��i��9�<�����eÙ`�exI�<-�V�M�6�i�*�OrȮ�/�k��ŕ�t�T�eo�f�Fᦑ�'%���.�p� ��+~