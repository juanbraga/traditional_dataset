BZh91AY&SY�7� �_�py���������`�z�Y����_GmH)JD LT���hГjhd�bb2C@�T��Tʞ�*@  h   �~jHbd��@�h  $ԂQ=@4� 4 h h @iP2~�1 L��b&���&A4�Q��~��O"SCF�� z��<�=B Zf�$0�XH��w�q$�4g��C��H�A��R'
V���WX��ݵ��e�b1@Q���f�������� ڊ��E���R[o$h�_R��_�SG��{|�hP��5�.ܪ|3�S.��r/m�L!��	�04;%	2f���{`�[�E%F^�آ՜V�M<Z���9HrkY0q�X��dጉ���4�V�+o��L�FQ݌�D�z��H39�;Ko��?��/� �b/����&r��6��PN%�;������QP��]-W7K��)�"�U1�<P����	�Z�ɧ��ϼ��4Y(�lkO���E��2.ﻏ��vT-�6kq����y�QƷ����.�����xu���$�YҺb��*Ļ�/@՛5�)�����V��qe���l�������HZ���r���3��U�hS�*uS�C�`��ph  
��L�(a$@��BH#&X�!�4���J�s-K��
�*t��@�����;ܳ��r��1���.�6�37g=�"�(Na I.����g�fP�1.΢�����Q�r�ϯN�e�7[Ě���{l��u��`��45f�cgx�mK�F��՚dN7Q�763�5�����j��]�?9	�aH���e�n1���f����4���@�AI�p�������6�m�Th0tNe�h�Sk*�Qk�7��)�j�f�N���.���$r��纜"���]s�ԎokO�r������?�����ls0'&�E3NT�hԅzc�\3��}���!�/eVb�}L��_� ��2+��A$ hK�n�۶`��d�l���~�m�2Z�ʲp2lZ�3I@0�$,�}Ba,�)����	&	CS�!��HӍ�ԓј�9<Ҁ@Z���r~�{�4�%UW��X�����T�^/� ������`�{9vW�l��>�ø�'�e��FaDi�r�5m��1�9 ��?�j�����O��ε�" �%:���ړ�-�{���9�Sgp����~�2 �Rr� t����v��+.b�2������*C0;�	�Ѻ�B�X�!S$�Q=p�m��q3ٽ��h:\�&�W��c�5� �X�&�L��G���I�d6)���� "X)֐�%�?*D�Y��aU<w�J�x�s$�w�W����A ��� ��blJ&��g~���oөc1X�4���`\8�3b��)ac�j��{eX�B ����m����aߒ�&�9.g\� �t"��=�3��J����0c{2���@Т��׀U$F�x�����}���(�+h�lI��&Zܦ!�6k+�̤H�������@�P�ۗ���S�4@(v�	�ӞU�m�9?�f��G�N
����3��jy�RD9����`�Hu��:!�� ��-:�X���Qޝu7�A�'$��`J)B*-aӑ�S�T6m��Ѫ*r����LuRƗ�f�E ��s	�6\�y"Ƅ���7�t���^/�cB|xb`���E-3\�Z-��ߧp��R��Y��:�X̸��s���HaN���c���"�(H ڛ� 