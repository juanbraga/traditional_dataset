BZh91AY&SYj�� 2߀Px����߰����P{awk��6*�DȏB
{�0�TƦ&OS�FF'�"���54�G����A�� �$DM4�OD�j4�ѐ@��`LM&L�LM2100	#M$�h���S��4��LM  4�bf��$O��]�T51\��!�Ӯ��@X��6�V����ޜ�~��i�J����"��1M�5�9�i�յ��q�F���9.� ��}��*�耕R��Q4��/6�Gm6�p�U��3�A��z�p�_FY��<k��A�)�׺D�A��6�\ʼYi�ģ�J� h��#M�i����îW���5ptcco��l�	�u=�tP�����&�Q�ܦmmU��屖�P��G�rť�C�1{
����0��6�[l�vʩ�*���9��l_�?ڰ�?�/n�~����p ����8�Z���d)��!L�o��e=�YpZh<>�5��k�w:���9Cu�� 6'/mb����Ѩ�j ����G��{i2g[F2�v�����3�vV,`�3
��Z�^�>�H+�9��r_��Ӳ��f�~]��2��"w��S	2gKQ�8L�3��a����g*V�c+����	�Z
¥2<�,C�sCp1E	��3�d�s�����\U'#�""<Z��4�H4���c.x(۩_z�
�-��1ʗ>#�mT��w�,�27���i8Ŕ��Ǿ-H(=��Xb�D'%-$@w���]z�@��H�'	�Y��Yk*Y�KJ������Z��*Ī��f~M�{F���7�<�!�������iXs�J��JN.����z�@�7��X�}�@7�E�n�6�Ari��ٗ��2�J(ݲk:*c-e~D��������d�y��c��Sd����:��gX��+��"Hi����0��dU�$�^3�����ba�(3�ņ�fYzH��P�ś���2��a�n]ykf]�E
t���Y��:N&A�x23vb�H�
�T��