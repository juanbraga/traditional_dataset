BZh91AY&SY��� �߀Py����߰����`��u�1̠&���JAOI���&�z�SM4    i�����      2d�L&F@��M#4i��ML�CG��jh  C���4�	��0#F�` A"�Mi��i�4zS�aM2 ��d���y�I
�U$�A 0A��J��>+� �ϕ�Ysm����5����B(�iv�l�
�,kכ{0{|�'D���m���"mM��I��Сν�T�t�����d+)���%{�o:�B��9biڞ0a!rB�1��Q���|1�U(�q�;�Ȱ�Plc�f7tR���Ra*FS�P$����!>y/+�}��lˑ�-���k'.�^|�@&���U�q.w���j�)�n)6p0�\4֮��^]K)Z������8-,�z/��r���;d]��L�`�D�s��	T�݅Bv)L�ό荛)��D!��2��[aj+*��΢p� 8�l��웦��)�=�m���$+1mi����S��˖��@`#�L��L'*��uq!rԎ�NaX!��DDMƅ��|�P�+v^���[K�ԁt˃W��/��җB�ɢ�����a�nm����@��O��z#��<<��(���ԝGT�c!�S _r6������26P��$Q11��J&gGa�!��K .��6�NJ�� eh�_���f��
挬�i��;nlŷO>�	QƆ�?���>�޽���Owo�������e*��0�M�<��H ��4;��ٯ��_�pn�0�4�N��
� ��ti8n���_�-/��/NKB����!�K��V��"Uu��+ALH`X4M�v��PڡX���@+;M�����lle�E�9�KX�I+���D&D���#����rJل���E����ex��;4"��7H��c��I&��cG3@I�SRN��k.��쨅@t�ˋɟ�T�8�S�*j��D�
�x��K�V�$<U�w���`V��ѱ)�j۩0�n��� ą�IN�n��zY�`T>&�}���ѯ��u��L�[5�ڪ6�|/�çt�ʳ[���_!΀F�6�z.q�xkM�=����v�u�w�z�1��9Z  �@/ػ�f�4���k��L.O�"�CĢ]�!ebhcE�	��w*dh ���ێۥ9����"�r&{�"�+ҵ*U���L "�P�,��(�"H�,6bl�rٞ��Ѐ\��%b]{�DX��PGa�~��|C5�Ȼ�0D�%�U��`�{�I$t��Ǖ*�c@'�w��C!�I�o��R\j�Cϸ�^Ӷ�0F)h+U��(Ɯ�2\����67!����s7��J^��%+a���,nTD���+
(��#� ����j�%����1j@آ�	�4�>\���W-��r�����3*���wg%Y���.*ΰZ��D�.��� ͪaD{N��X�ooQ�d��0VGrĐC�]��BC�Cp