BZh91AY&SY��d� �_�px���������P�8� ;�j��(D К&i��L��)���S4�4z&jz�S��� M  ��  JbQOM)���0� � &�2d�b`ɂd ф``(OD�S�?S�<�O(S�m@24�54H�
�	bD@@X�D���. �wuL����A��~���H�`ch�d�Z	�[٨׿�B6EO(�����h�k,D����D�wB7�QX��mƍ��n�r]��!BHcj*-sk���铤��kղ-�֌��܅u����-Tb!*o�BJ�wL6c��ϱÄ�!�2f|���Z[��_9C4��n�/�]�߈���!�w�������h�([O�Xˁ���8�P$ׇ`"A�P#����1��Jf��r�h���Y馀�e�V`��`I
a!�"�An�n�7��ֲ���J�0B��|�BҘ�B��6�ʑ:e2��	Td�E8H.�a�e`Z�XMJ�1i-&)KoqX�,M4%+�"�!SYHVV>�2�����U�m-ar��h3�I�v�#S5KUk�lnԋu�Ǭ��
��v�2�м��q�b���3>!��:�n�Q��6���[
s�8G���?���66����!�d{/У�%y7�"�n��y*9U\�2a�L��T$q���p(�Q̃ Ma���(e.��b0	�-���O���Q9�p��]�;��������y|?�be��ˆ��OH!��}��΄"��g��A�>���e�?A�Yx�7 $#�W~��W�ս47�ĭ;�B��!�J��*�V'��kΈ��gV`�}��yd%��"�kg�=��&T+��-��6���V����{)��9'��n�7մ��B�����DyA��d��H��C�L��k�6*98Bh�XP��C�j�hP'� `ޕ2�vXc���\E�0!D��T	�ϕ0�_B%$�1�:�[��Sъ���S�0},)�VD�%qZ;I\�S�;���}�B&hfd�_^���Ҩ�a)bR�p��I$1�!�Y�V�[�8���B��-���Q �F��*İ�m%s��]0����{]>�CMlV)<`"]0�����!D���tm���Q��B9A�(���C�I�<��0纫ӊ�.k�q���6��MF갱U&_ B!��	jL���fW��!���EE'���h��řT�/D�eX�~����hEA�;�5�=}*��YM���(�EŒs�C<��Q���!`�;����8ˑs'	�iJ��%s�g׮v[-��bqo��g@�[<�]�oxҮ<[T�٩��B33/��J��T�,��&A��;����"�(H`g2n 