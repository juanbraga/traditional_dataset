BZh91AY&SYSj� �߀Px���g߰����P�Թwv
�XIM(������A�C@4 4��S����6�h�	��HH���COQ��'�P   z hsLL�4a0LM0	�C`F"���#!��Sѩ�ɠ4 h�h��! W 1B"I�{���f��Bd�?Rp�$�"l\쓋mt��=Z����}je{���Q��&�hm��7G22�z��ͬ��"%F3!(WH����gqXde�d �J 
���j��v���&4��;qr-ry��Ý-�ᵨ�n�C�����"pr�+YЅLϡJ����
�����!A0��&��%$9��4�2�F�vIQ�YNh�V������m�lm�m�I���{�lFݤ�V,��z�ݹN��瘺W�Bf.Δ���9�Y8�u���y��llr��٦���;��BJ%�Vt��D�>�s�Sd�)гwS�	P��q���lF�-�/)ҩU��E����#���-I�`ơ9~T�
��i���gһFjB�x[����&�hbʎ��0$��h9YY���M���`�EP��0Z)]�5C��$�CV�k�*��qE�]��si)hF��"�'
*-!0�����S�03e�(H �X�s��reL<M�B�اP��y3�ڰ�D¤�ؠ����VfQ:H�c-�)�U}fQ
��cؼ.T�Z��L,0� ,���b�����V�[C!Dh&�Q�)^�Ւ�XÉi�����R���d�j$�M��F#&��΂�J�2e�:�7;f��!d-�@<}��5�˂7�D�F���6�8�KcB�7&5��r�,�1�T�%����*mPP5�E�@u�a*����O� R!KMWU�dj	(�d��hN��@�0�ihZ5f&Sň7O$]v"bp��A?�q�&��"J��,���,	L潇]_�F��Z����"�(H)�|�