BZh91AY&SY��� ._�Px����߰����P�s��w�H��I"h�j�h5S�=S��e7�5SL���A4ҕ0 �L     JdD�҇�24��dP  OP`�1 �&	�!��L��Q�ԙ�)�Ѧ� �i��(���%����*^��u�/j���H�
_���']ABPmE)QF'[��զ��,m^fuDNTR��Nf�q���K��[��%�":A1؞�tῼ������N� �� �	�LS)�^/�в�E����0���)�tB���p�_i+:����4$!��Xv�7i�ű��
浭[RmjZ���q��@(D�N���z��h����쐹�01����w
���i|b;�*���T>�U@�Q�� 	�p�a��q��b����k�zI����F���� �$kS����٭�VΪ�n["�ˣ'3q@�[þ�In�jwL$���Lky�0�:r��e���C#�O�`o1�R\��d�������ӌ�![35S���90S��0��p�ow6�-�vs`�jc:g�"!��<�Ii��b�Ɔu�N"!�t����m	��7�iN�{�aE�lZ��/,N�f*&���]T�Ȇ̫���32�l��cnv�	�$$$�i PDb'����I�oh�nXs�u7E.�ɖ
[�D�$5%D� ��(�
)3��)b%&ʌ=�ى�c���m�0�J�t����w{U�F�ϫ�i�o��㇗��y�>?K�ʇ�;���㿅{	$��v���WbQp�[���6�1y�̊�GO_:�}���/Z.rk��1��oH�P똄���7�NX��i�*��%ǚB��W7�A�z�C�j�?\�����"�%?l�K9�U�����*�U6>wG��,
g�-0���=���� _�r8�f��pq�%/�
@x��X+h�Ք�ԛ�'b0�����
�RHR!ַ�^N!����5P-f\
9�k�U���4�L�׳���YH�Fҳ"T,{K]�pӶ����$ Lř�|����Q��{�J�8�9Xp{��f
�eu^rm�
�����`Q��p
�����"$��~����~�	�X��e޲�_b��!K���tDȠn��:��e��A�H\�Cv�p��}���>��0�i�����h�V�'ћ,��T���誜D�8M�h8$_| vΡ���j5tJ�E,2�f�3�Ok��3[��-^���=�)�Ѩt
d�~�x��2�ŁB���B#;9�``�0�M�
���	Nf9�:�~6L�hp�0J��jG��ifp��M�H�Y9�rq��V�/q�B�>U��92\�2Z[��F��]��BC�WK�