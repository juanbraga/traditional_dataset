BZh91AY&SY'LB�A߀Py���������`ro �  ��Q@�            Gt�   � � ��       Q   E@  ��  @ 6   ` P�a  B �    B !  �    Q  �P �  �N� @ �(�4 	��hi�1�i�<S'��= �M���R�骞�        q�&�a22bh�A�L 4�IEU    ��F0RQH�Hd4i�M  � � ѠT�j�Jh�42���&�� �&�4��a��p�3E��@Q�]�
�(Q>R>%�H��s�������|����m2O:�\�Ư��m���RD�`����(y�f-c_g�v�����|^ϰ�������V�lM�lKeV�x��0�w�0�!�&�[�R�w;�M���b���l�w�N�)̒��`N�Nd�19��el��-�\��6Il-��U�-�)6U.�`�6���Q���l��$���0'�T5GGW�)�.<i�g�m�sľKflP �3@)�� E�� +h �� E�<� �B2e�'$�bg�� 6Z  Yh �n13Й��;����à�h e� �� Z  .( e� ��dD� DI�dD�dȌ�6˓@ �� �@ -���j���+�q�����[l �����p   8��E`  `  `  `  ` QF r(Y@l�I�dD���bL��"&aM  `  `  p�  0  0  0  0  0  0  0   "I��I�           �  `  �� wt  ��  7w@ �� wt  ��  &�  8��           	�� N6$ȉ22o	��s&Lɤ̚L·�uQ�HA�13=�'��13'6�m��G�lbf�n1=\�,I�e�L�{ ��h e� �� Z  Yh e� �� Z  %�  Yh e� �� Z  Yh e� �� ��  om� 7n� �� �� ��  n� �� �� ��  n�f���������xNs��8Ns���3134�|q�'9���M��i6��l�S!2v�8��  ����Ě2@���#�K�n�M�@ ��  �fd��I3�37,I�L�&DI�dD�$���Ѷo$���;bf&a�\b������ Z  Yh e�n� ��n�IbL��"&��c13134���DI�� ��I�͠GH�K@I�9ɝtK@ -��ܲdD�d�$ȉ� v6Z �-  ,�  ��'g�[��*Www.y�Y��9�'6Y�څbb��A1��d>�����R��^��B�m���a�sQ"�$����(l,F�� N׶  �I �K��I~I$�I$�I$�I$�I$�I/$��:� �I$�%�I$�I$�I$�I$�I$�%�pI$�BI$�I$�I$�O^�@ I%~I�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�K/I$����{m�{��{��I$�I$�I$�I$�I$�I$�I$�I/$��I$�I$�I$���{`         ��  �                             ��                                �`     @        �l    �w�wp     wp��             ;� m�                                {�����  ��I$�I$�I$�I$�I$�@w]$�I$�I$�I$�I$�O�I$�I$�I$�HkZ�I$�O{�I$�I$�   �I$�I$�I	$�I$�I%��$�I$�I$�I$�I$��` I$�I$�K�� ��l � �I$�ǽ�v��I$�I$�I$�I$$�I$�I$�I$�I$���I  m�    �I$��$�I$�I$�I'�$�I$�I$�I$�Iwp�I!$��� wp �                ��          m�@� �                ��           � ��$�I$�I$�I$��	$�I$�I$�I$����� ;�   �� �`   Z�I$�I$�$�I$�I$�@Z�I$�I$ �I$�I$���K�K�  �I$�I$�I$�I$�I$�I>I$�I$�I$�I$�I$�I$��$��I>I$�ִ�I:���I%���I.K�v��I>I$�Kϒ�I%���I.K��G�i$��I$�$�ַ�.��bI)$�I%$�I-/I$�]%�I$�$��II$�I>�I$����I.���Ie�$�K��$�^Ii$��I"I%���$�N뤀��  m��� ֵ�$�I�ll�l1�<�[�Tڛ�i�
	��5UT@Ʒ2:���;�~?C���AH� b!���O��د�����)Φ"S)�{�2jj7�%�[m��12Hə�L���2"d�Y�2fLə3&d̙�2s�V,��sG3'8�fLə3&d̙�2f�13131ݫ���2fL��8����IԦb,ԍ;U1�D	��I�<Դ11c���+KL���w��ke�[�s1P��JS�ZִD��I$�H�$���Z֒I$�I$�����I$�I$��� x  �� w      l�� -�����        ��qt�I'�I$�]t���^�Gw	%�I-�i$�K�ۺķw�I%�]$�>�=z�֒뮒HJ^��m�  l v�v�`  6� �ۮ�Iw]$��m���	%$�mi{�u��y���I$I$�^���ׯ�K�����]kO�I$���$�It�I/Io��$�ם�כm���J��=��w�o����W�~_��K�˽%�}�Km�1���{�m���� ��]v��^���]�cm��m��G��^�t��%�륭yj��\�eS)�M)4�%_Rַ�|�o!O�%��k<��Yv��J8�mF�LG�mFҷ>D)q��T��"�	Z����)��S�����3��jy��jm�(�Dc�m�R�#ʧ��[K�-�>������R�"nfgR��hZTלI�^y��C��R_<��{���ϔ�6�6��|Sg��cНO�L�a	�U�Z�ZT��zq��-Ž�K�y�Y井�e%�)(q�ͼ��-�DyM�-�o�Ty(G�*QWp��K]�J���Z��n]S�8�iS��o�<�Z���<�,�K�{qJZ��[�_��w�%k�H��'wxc�����{{�ݛl���ҽ-w޼֖�{���]��=�/��]+[K��u�k�t�&�nۭ?���ww�t�%�u�-�%/1��y�%弃ͤ��n��V�[�x��%.�u:���L�H���.)6�-kQ�B��~[�R�q�yiK����S�RV�ǜp�_J<���V��<�RP�)Q)��եk�Zҥ8�n)p۩q�m*|�|�[8�yn"b<�[iv���<▕:�iR���u1SU*U�n�gR��h�J�p��u�oKn<�ި�y�∮�ϒ��m��	Z�!��)OB�?=UJ���j��F�kB�kN��B�|��R�-/TDq�m�V���Q�θW��LD��J|�>�]D%�ժ�Jֵ�h����wl���]����u���^�Kn��[ݯ]/p ����~ߗ����[Z]u�Z�{�+��^��~I���|���-iR�un<��m��m�iq՛c�Qo�#�6�i[����z����w˩���R�u3:��kBҢ��R��ͼm-�Sk}qy:����R_!�[R�[my���5Z����L!JU�Z5+Z�,��q��U>yHCe%>��"�bŌd���&��0�4�Qə3&d̙�2l��#��v�k���)�CT�#��!�5��k����S�k�qѦ��	Ahx��҄t�J*�.���kR[kΧG�<�H��ml���Z��d���,�F��8��B@�Dc�,�CT�6�5�q��!�5�C\C_����7{v�k/sww�t�]׵m�4qk�RAh}�6�� �8�k�hjq�68����)}���R��F�A�>CN��|ۅ�� �(��{���~��������^��v{�� ��o=�{l���t�z�۷^�^�]���k�wr���)���뮒ֳ�%���u�k[����u��ZVڶ$K�C]ZZ����7!��H��}ə�-�i�C�H�C�j�|8����kU��b��]C�k�k�mPm���ZP��T��"�	Z���M��>A�� �!�6�����:���K��8��!�C]Ch=q��CZ�)q��	��b�q��֑hjH���غ����*�7S3�Jֵ�*u�kV@���W�mL6�bN!�ZF�����!f�v5�4Z��q�lm����������:����6��5�B�Z��}�ze:�*QWHJ-v��f���(:�!��+���b�1#�kTCX��1T���j���m��[�E��HCjߪZm�����c�5���!�?�r*Q�E\E���-iR��X��k�k��O8���F�Ah|�(-
m�ŵ��uC)��^��khsik�5�8��c�Y�>CM����4n��3��R���+D\UM_�m�y���������^�-v�뮗}鷘ol�t�{�ϵݥ�Z����/�������Л��۵��o{�Jք���h��j��^bvq��5����mu��F1qhk\B�ZC7�)ch)C]ZE��OQl6)kd5HRǐ�ɉze:�*QWHJ-v��f��)uCN��qbB�5�
 Mvfq+֭�D���5ť�m��5�k�����1:�h:���P%��5��"��J�U�\!+]��	R�����)j�#�(����q|��qз>G�i�|����P��2�)�kdCV�D�#�c�[^u-m��!���[׋���Tҭ��ԥkZЕ6uj���KCh���8���-#�KP�G�#�mj�k�R�ˈ��-� �6��!�iz����Y� p�Hj��<��!�*QWv�"���K88��#Z������1�[X��CZ�)o�U,�<�(8��k�H���-�bG֨���p�hk�� �!��Q���ֶ�4i�w�~#�Bԩ]R����k$�{n��I$�kZI-m��I$�I$�S�ZI$�I$�N���  ��  �  =�   ��� m�wn� <1m� m�l ��   �?  ���z֒I:뤒K�z�&��^���$���-�i$�	%��v�ğ$�뮒O���c޺뤖ִ��[�x��     =���     �kZ]�$�k;� $��6ֽ�]t���^�I%�kI$�mukפ���[K��%��攒I$��$���$���wz�� ����s|ֿ����m�kZR��j������c����m���l.�]ں���֝u�oy�3�;^�/Z�KJK�I�-H�&օj!0��Je6R�q��v�Z[ZJ�iZR4W�f'��,qqĉZF��7�x���ub�6�hb�LKZ�A�C%��S���F��<�Hmi�]LT���h��F�kR�*m�գ[C_!�����,�CLC�-!�TF1g,��5M�MDc�z>C[ZZ���!���u�k]B�ZC7C5N�5jT��.��Rֵ)f�ZCX��F���b��5�!�B�e�c����m��i�6���r�Ck�֨�i�#�8m��"]H������T��])R���ZV�E!jCiCX���Z�o��[�:�:�%��5M�aKCPĊCZ�x�+M��:������u��8�)����6���&����b�U4�DJөJֽZ%M����|�+H����R�!�5_%��H=q��CZ�)Z@���)g�mi�����c���!�!Hj���_���{�KK��%������wp�w{���m�{tK��W]eݾ׻��w��g�+R��D�B�l�)�fִ�V�^k�{�>�׾Z�g��]{I*R�>A��hu?�AMD~?�V��B!�{�Ȋ�lm��������8���n��!�!�Z��<�͡���b��=��R��t�J*�5iZ����H���_�g���k�u�6�PҜm��B�T����(��5���+H����)mbC\CX��-���J�T��U���+Z�J�5�:��- JB�y����uC)�b���jѪB��JA届Y�#�i�:��$����q�CT���y�OB5jT��.��R�IMpb���!�5�55�B�@��������ޛR�R�K�aM�R����0Ķ�:��9*�W�)*��ZT�B�-H1�%*�#�ڇuť��!�1լ�7�N��\u+u�bq
q�jR���
M-e!kZ�d�m��6�����wvm�
Z�Meuֽ�u�K�^������r��i%ҵ�).���Z��:kkn�^�ե)Z֩��Z���6�js���>tũ�,l������)�V�:�.1�mŶګ^B~�=2�Z�*��B�K�D��S�6��\D����[���6�)n�mg��l:뤩Ly�0�]q��o�v*U)�jD��5IR�*Cu�mߢ8�KΥ��(T��b�r��8�����),���Ej#�z\>~>|��y�X�����!R����t�UM)d�)Jִ\�M(㮸���7�0�y�X�5lV☭8�m����K�n6yJBV��[n��s^BkP��ujT��%E/T�.c帳�z�1�=g[�KS�>mo�m��u�]tꖷ�[l:��e����_��|��I,�%�=�gwl���=��l��Z�֝z�-�����ߗ��z��6��Ӽ����u�KkK��KZ�˗[�g���׺�{�u�
��!n�R����O�Z�|뭸���C�9e>�y�Kbu��,c�C�[�Yz�oҺU*���V��+Zb�&��]mԭķ�1p�T1k|�c�i�>|��u�b�:�[1jO�ڛ6�:���Lס5�ze:�R�W(Z)z���\m�:�|�S���i��b�|�8�6�T�Y�)o�-�b�|��J|�L�v.�W�RUq��v�DZ���%JW��UK[���mN��q�ԧ�<�l|�u��jclA�8����WJ�TҖM�P��i���J���:��\S���qO��1Gu�-n<�1Jc���mm��Ӈqo�Jۈ���Ze+Z�Z"⫳�6����{o{;����u�׮M�ֺ[��F��`v�gw'��)KkK��KZ�y��[�;����Y�u�{IIQ�:�V��-�����yLb�y�n���)�9�6▗_,�b��n'�nf�軵^�IU�jҥ�jvP�N�h��#�R�R�K�x��)J|��b[u��m�� �\Q)�������SJYu(JV���)*y��ť��C�1�Z	�7�N��\u��J���ԥdGX��8���oT�J�=իU*��B�K*QG�|ꡉS*"Xٵ��-o-�Sέ�U�RK�q��qm����1�uf��3U�]گT���5iR�
��:�ΩM�qڜ|�����|��8�*SϞq���-޸�܈�!�κZ�?������*�����JͩKT)Y�&��� )��j)(J��߿�����C��{�w�I$�ބ���I5�i$�!$�I$�I$�^�{ޒ�I$�I$�� ��  ;�  wp     ����p w�.��`m��         msgI$�z��Iu�I-k^�i�I%��]u�I>	/x�hI���N��$����ϖ��%�]$��Gw      ���m�    w�f��%���M�� 5�jI����뤟;�^��IkZ�I%�k��z����ִ��I-kbI$��I$��k��%�;��o{����������{���o�Iw]$I{�m��l�m�z�m�z�t�Y�t��eֺ�}鷘ol�t�{�ϵݧ��.��KZ=�.�ֹ�mm����׮�K޸�U%�X����-��q�8�y�7�����8����ڑ\ɉ��!km��y�K�jժ�\D�h��(����mlSt��Ĝm�8��ib�m�ϔ�%ll���\q(S1�8��{�nf�軵^�IU�jҥ.�-N��m	c㏛[��q��x뮝R���m�\[�R�e�c��
S�=���T��Q��kL\DҘ����[q��ּ�%�#�8[�:����5�qk3DN)�]mԭ��	)թR���-���,�ώ�O/�1Zu�\cn�ť�u��bԟ��6mjur��.��۬u�JyO��K��Ie޺^��l����6���cm���K[u�N��K���������n"QIZ�ZUI�-H�&օwu�~wm��g��Y�|��[�-~�S��SQ��R��u.<�8R����u�m�6�&#Ckl�)�F#����%eTF�+Z"�)T��m����S��yn8Z���-���R�h�b8�L��g㏜u�n�����ve:�*Uq��z���M���c�����[�1�\ckn�&�8�|�V��F㮘�=,��~�k��^�=�֒�Z�m���)ן9�[:��:�m�-.���1�cm����!ŸqK[�G���e5IYU(JWhE�R��][o���)��Sm��>|�ǌJ��>q�� ��JU،J�!�qi�<��V�L�$�z�k����w ��{�;��`����Ywo���w��`��G��{�u��Ȼ���w.�����Ӻ�Z�*���-KԥD:�Z�cx���u�R�R�1
q�jSב*�8㏛q�9�0���1j�bW3UȺMjԉU�j���
Z�8����届y�ۮ��K�q��qm����1�uem��:�~���u��P�r�	�-0��JR���)Ju����y�[8�%
�3`\�4��;�;�KKM�6��@b�XP$�9� �y�b��q���?]�P�󮖥����q�wm����=2�Z�����-K��M~��TK�1��c���:����M�\��⍸�Z�S}F�]c[1+���]گT�E\F�QkZ�֝:�m����K�n6yJBV�ϭ�8�P����,�ި�c�6�uJL1�-Z��&�xc���ow��s��w���Z�Meuֽ�u�K�{���������{�u�).���Z�ק�'��u�w���JT�\E)N��ky��yn�뮝R֯<ژuŸ�-f\F18�JSٸ��<����[U���E�e+RW34��iJT�>uD�H�8[K��>Z[c�C�[����'�Cn�ouN<t���̙��]�^�
U�j��	��Zu�\y�[b��:�[1jO�ڛ6�:�Z�Xc���c����8�jqm��ֆj9k���Ҕ���h��R�yjuf�%�8��)K|�m�u���X�Ș�b[d��ٸ�U-n6��m�<�oGQ	�!Us3HZ���F-�KR�c-���RV�؃mF_�3�q��:��\S���qJ��9
f���kZ�Z�f*�;��`�s��Ͷ ���k��O�%�t�r����p�^N���׭JKZ�u�%��iiݳ�>׭g�����j��N�|��[�1�\ckmO���[�ҵ7�0�t���Ko6���3Q�\L&�jJT�JT�-JS�>m՜[�8�5qf�Siu��8�-��q5�C�p▷�#S��VꖳAoG2��
���BԴ�*)�
R��1՘���>u�\F؃qD��8��C�:���l!�1լ���&{w1wuz�R�#P��hZԲ�u�R�R�1
q�jSב*�8㏛q�9�0���1jb��ͭo!kc��V�k���-IJ�)J���Jyո�ζK�q��qm����1�ufޘ�c|B�)M�qީ��[��Yi���*䁚�
�F�c*IKF:���ߒI$�Om�$�I$��$��)$�I$�I$��֒I$�I$��  �   �� ��     ��{��ضͰ��� s`     �����Z�Iu�I.��$ֵ�i;�I/zImkI$�I.�;�v%����뮒O��lz��]%�]$���{�x     wm�f�    �{m�$��I$�wm����I�t��뤓���i$�ֵ��^���zκ�/u묽$�%�[�)$�I,�I-kZI%��^��u����}}__��~{���%�u�I%�=�g�m�{�����m�w�t��k�&���ݯZ\`m�;]3������]%�g����<���k���ץ�]�u��ۄ�Oǟ�0�]q~m�{q�;�u�Կ�6��q�[o�q�q�.�zg�swW�E*�5Zօ�K-�8�;qO1�!������̘�Q�q[jo��ckb��'N8�lm-��b+���M�Ԕ���hZ���u��R�6]��Q�Ԏ���KVq/�q�m�6���)�6�Ͷ�5H�^�&�!Us3v�*҅(�n�R���m�\[�R�e�c��=��EU+�[��ִ֝m�͸�:�WϞrf��.�T�\F�KZ֕�e���K�qq�qk3DN)�]mԭĶ��8�S���:�<۩�z4')c�Z֙Jֵ�h����x�`�m�Xm�W��K5�{�˭u���o0.��z뷼�>�v�����]%�g���^���ik��^뮴d�����6bԟ#jl����%׌q���[z�1N8Z�[m��1�q����F��m0��
�����S�)N���R�ym��i���q�1ő1�6��R�\F1L�n��n�ڟ6�q��?[��u��������޴�],���.��-���8⌿�g㏜u��Z���8�p����#M��hZ�w���mq��Z��RP�-R���>q���<�-žm*S#�8맔��ŶR[yֆ���c��ͣ�qLb5�G�Z�����JQKB�T�E-O�Yǘ�-��#�8�=Q�6�Kuj-հ�d�F��=�i��kU�%������x���m�;��6����K[u�N��K��������Ӟ�^�K/Iu�޴��z佽�k_��w��1�kY�}��E�)*Y���-��!������%�u�%n���c�n6����#���n���IBT��JC����"<�6�Zi����K��c�b��%���[�[�c�q�c��UJjB��f�)E-R�)n-n�>aǵ�����mD�kF���Z����V��kMheyN��:�>b�b�}�[�q*S�|��]�]�ܩJ��եKZ��,ۮ<���cî�v#�<���Ŷ�m����kZ��<�ۮy�lF9k���-IJ���kR��1�Uܘ�Sn8��W�x�8�>b�ӎ6Ÿ�-,S�,�Q�<�]�fIn}��w<1���ww�������Mk��u�]ڽkޗw��g�7�t{�"�J�[[6��k�OZ�]{���ȵ!Us3v����B��N>Zҏ���b��ި�c�m�6���)��S��c�J�������]�ܦ�Ws:��kRV��b�u��ʈ���Zֈ�ʥ=��EU>Z�qŶ�l1���y�by�>o�Z�UKRR��*Zԥ!�:�+��m��|���p��NC���:�o-�)�)�:�1i<�m��P�RW37iJ)z�R�qj|�%o�y�:�R�7+l��Zި�b�|��4�Kn�LmFҧ�霻������*�5IZ֤J�gX��-�LF1���L��b���SkK�aN�;�|�8�[Zk~Ķ�aKU���|�m��;���/y��wv��{��Y]u�w�y�����kkǽ�^�]kJK�뮖�n]ב[ijR��*Zm��L��gۭ�덥��C�1�bu�]q
q�1�SmO>F��1(E�
������DD�Ӯ���Z��0�F��伖1��y���1O:�qo��Sn)oW�yS;�������*�5IZ�B�q�)�m>��c�Jި�Z�|���Z����|������6�޼�|�F;k��U-IJiHR����!��RU�E�I|��mI[�c�!�l�6��k�c��-/}F��bP�RW37Zik��R�8�嶖�Fy�1jb���Z�B�S��[�(��e-խ��k]h֣F���7����Zֵ�d��zd�I$�Z�I$�I$�I$�K�{�����I$���^� ��  ;�  wp     ����p ��m�`�         ���.�I$�I$�뤚ֽz�wp�Kפ�뤒|$�w۰��zI']t�{π�뤗]t�B}�     �/l     ��kZKmi%�I���  I>I���뮒|�=zZI%�kI$�]��ׯ^�����o�H�$�ݢ�$�^�ZI-kZI�[N�z�{��Ԫ���5�i�y���N�YHZ֫B���۳�����{{�ݛl��k]/i�������k׫�v����ǽ�]+}�H���%Uq�{m�3wsuw:�E\F�+Z��~��o�#�m4mJz�1�q��|�qÎ8�)��8�n��[�y�e�*�jJ�WhR����!m��v#���|��|����s�<�1�^u���І)�<���ġR��f�M-s33Jq�[B�J�F�S�/�8�jֵ�}�u�--��y.�ll��Z�u��]�]���iq��k"�F:���ި�c�m�6���)��mo�q�8�ÊN���>[l8Ÿ�j-��.S4�.Q7z��i��Rp�jS���yUO-o�qm���\RR��-��qIy�C�q:�G�����~N�u�I%�=�gwl���]����u��:��ooz�-���� �`v��{���֥-�.��-k=��i�ׯ+[;�z��\�{ڕ�m��q-�a�K�c�8�o���c�m�R~Fԭ��ݽik��oݻ��k��}��^�뎼����X-/�kz�1�q��Q�R�Q����8u�>b�m*�.S4���3WZ��i��R[�R�q�-ź�֗V�K�ZJ_:��|�ul�[ci<�}�"�U\��!+R�w34�6��O[m����1�bu�]q
q�1�Sx�ԝj�:�Y��m���˩������M"�#T��ȴQ��y/LF1��y���1O;�q��N1�6▗_,��-��fB��Դ�V�Z^��v{�� ��o9�q��;���Iפ�o���.��o0.�����r���Ҵ���뤵���޽4[z�g���-7JuөE�1�6�Kuo�0���k%/>y�Ko:��q�1���z:�"�����BV���%JI��Rz�8q��<�͖��yn��18ojVDu�6�o����멫�����M"��u)]��E1:�)�Kmky
yLb�qn}�kF��F�""kZ��n9+Hm�)n*������TmoCӫ�L�P�Rj�)R��)N(�T�2�%�u���}�[8�T��<����qo\F16J]�cщB-HU\��!+R�q�1��yŶ��.Ktu�t�u���1�!�mJ�L�)�m
m��i{�Z�)Z�wt�[=�����m�{{�m�{�]t��]d�W�.���{���޺g�����]k���֖��r{����׬���ԥkYQLu�'�1�ӎ6��[�)�y.�ll��ZҎ�q�c�Nއ�U,�L�4���R���R��8�D�c����uN<�q*|�Ka�-�-D���Cm��Ρ��%�!J���%j^��&��������y���y�by�'^c�I��#���|�S�컘����)5s3�Jֲ���K�1�Q�|�S�_c�ڒ�jm����Z�|َ1�"��&urɔ�JM\E!j\�)M���[�c�帣n���Q�)o�o��X��-�LF1���LȆ<�ֻ�뤖��-��ws��M����`$ֺ�u�]��֝�]��g�v��=�\���k{֟k]r^��u�oZP�R�qJԵ�D�M���mi|��R��Ϟ1���[)��L���%�[q�mO�xw�v�k���뤕�i�����o�q����-�)��R��6�_�|�p�|�֦�G��|�E2e���&S0�Rj�)R��)N�ͭ�1�yո�o奎)��[i|��cŶ�Dcp�V�P���Z�(���BV���"T�R�-E����K�_6�m���\F1u�%��F�I|��F�K������v�i���u�K��WX�Hc�lmǖ�^cㅥ9�(�m����Q�X��?��=����m�5���6��a$N$������V�`���&��d �W���U�s.0R
�������ԥ�Ry➘ܔ�.j���Gp��J\ԥ�[��8�T�i�C��.UKϼ��A�¥㼒'��T�ܡQ�Q�*؇���
2�@
BP_����}�5H�`8$�0��tB��&�LcI������p�?(|�\��]0�?�)~Ou�r|h�����A�_��r�}����IO��N�������{�κ�B2��*_��x�|���T��A\���?�|��i<�`]D�	샟t���{�D(p|Q� (	�X\�HaPD���O@���N�~��%־@KPÎD�?@��N>��ATߥ �T����H�kJR��JP�|f�>�AM���ϱ3?Ǧ���0&',4�N�۬hǫ�!j����� ����F�#�S*��SN8k�����6B�O�:c+5!!�1�o���o��n��[�6��B��ʗ�^钓�H����,��Jbh����)��MP�MSYL�5LUX�UMMS�bX�I�Ȭ�SJ�S*���MI�Қ�+#Taa��p�����&�U���\>齳OA�:�.@��V)����X���'C�WT���qN'j�q�-��.'�̯��t�?�������~nf�} DA,�3(1@8�i�wߘ����<�&t�_� (&�Ɉ�������'xz��0�t����L�<�2��&�WC
D��?]��W)Oe5��9O\��3�}7�{\�h���T���Q'��@��8��0|�2�#Ts#��&΃ ;����PP��wDA&@Ђva�tB��% �bX[=��
 xB�Ќc&�2{�Y躅��8Dٽ
Đ�h
]&�;�pк�$��%�����9�\�NAOG�p���Xօ�-���t~ޟ�Z�݉�>�x �y��I�Q��t��0����;Ow�a�^3TH���R������l�zÀ"UA%�����{}�\�'�r�]���8Py�av�������(X!b�Uư���zm�2��i($��.&���a����]���Z!ǅ.�"	�nc�-VxF��be"WL��g�Jh��&�-Ӽ��{�,J`u��=ۍi��@O�����^ =�d������0x�N"����J��y��Y=��$����w����H���@�aC�s�ϸ4��w$S�	t�*0