BZh91AY&SY�'�� �߀Px����߰����Py�n�3����.�A$���	��ɦ��i=L��=!�F�h�4�4�#S�=C@ 2  "�@��2� @�Ѧ�49�#� �&���0F&D!'��OBz&C@�    $Hϰ�B$@�$(B|��qQ�bF䁘5��Ӄ��c�F�S��ء�׋��1�1���B���$5���wR���y�Uu��om�)�|�JI�j�?�?�xWV$X�.?J�[0�݌`���&D��$��D�:"&a�p_�Z֫LZ�j�㓃KHo�;��w��:�݄R�����<l�m�Cct����*XP�@�|a`��h���"0y��o�X;�X���Q��m&��"�Rs
D��$WʏEU��kxeA�U�r������uew��f�NkO6�!��66�Ͱ`�'�f�:�-�
&�eTݔ��&`.����[�J\41�s��Z!����Ng�f�j�M]Q�FV�b�;���'Yg��u�ΘwV�8�����I1���zq��
t~�����p�\��z��$�\O>��n.&+2�e���b���[�7>{�,Q����!��p�666��D�?�9�l�	�I����Aa�~�ǜp��+qF�䴤03�T�eÿ��5�����8w�!�.���	#��ݵ��Y�a�>�5B��͞��8L�5ȓ&Ί�	<ëP[�n�b��>�	B��V7�.!�郜��5L=\����n2]{U"��(N�&n�"��UU�0���q������ڈ5��(�U_�~�������2`䃂MZA��l��K!1������z���E*�"��P%�B��`.�IA|%8L���j�8�yL�Px��x�!���M핀�j���A�H1�,.
G{�'�?�c@z�c�j�[��5�FI�MF������5�i �c2�����I�Z���JQa�Bz��2�}y�A�H�Of���5�W.�D�D���$��yldY�9k�BL�k$@�$]��dhh�.�e�mc^�־Rf��!��"U�#�T���0r���d̨Y���68ᦦe�Z���r��K��%�O�
4�ܑN$.��|@