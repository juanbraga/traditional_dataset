BZh91AY&SY�8�/ �߀Px����߰����P�8ݒ��Ud�%!$�4i1h��G�ʞ)���!�1��	$L �	� � � Jd�i4H�j�i� @4�`�1 �&	�!��L��Ji=F���G�z��d�@���I����[�%A�^�Fu�X��sXb�� X���i@� `AP�9 R!�8�A��e� ��,�!�FJ���u-��h{�9!����ɹ��F��Q�ZJ�Q2�������ꄈ��6!>d��M�M��g����@j�DV��D$Z�
îZ������L�̚���;����C�ކ�O.x���������'>��5�FA��8��R#4Nz_��(p��YNFw����`$X��5��Jk�JԀ����+1�-�KA^���F�bGAeGVvbVvRv�1!�2���������Q	�q�M)�fY)ʹS:8�p�4�̋P{P;�ܨH�w���e*��
�(*5�9Ō���D$�x��#�y	d�vZ*��+�d;���wؾ4�X�L�@������S2�Lh�|Ry�fԐ���$��O/_�OX�6�vJ�/Y6������BQs)��JA|B��Z��a|	r����n�; �9Z�Le��$%F��.�gWy:����wzNr��:;�g���_V?���Ӳ�λ�S��ĀK٫��]/@��W��K�Qˇ��1 5g_+~WNB^bA&�pe�xr�9���*�%�tI W��d����iɸ�\�%yG��c��	��z�fY���N�Z�\�$�ݍ6���G=zn��c,I��m���'�S��N{M�yi�-�Z(w���*&�
�	A!@B��*�gFS��$�+j���Q�Q���B[�LL�a���tA?]�\_d���X�����r�����$���(��xHq�9FhҮ����e�G:ѡ�4�eBb:c���m�ټ����_�_V�#q�*la�0�M�����!��|�]��as��Or�	x}� �����^�i�*����wK&;6+�HB%	��.,YS*����YJ��+˘�n�p=���F
�ӬZa@p>I�c&��	9�����6�r6#�.�¤�鰉�(��|��ҽA�L���J��ٖ��;~�$���o�MF�ǟ,v�f}�u���j8��Po�F�Q�橰�U��q���P9TR�&q;��� �j=����|	���<)�L��(:4R\a}A"&�ܰ� �ffk��aCp�Ɂ�	�]��52]�
��Iq�6�������K=g���
���r7^o����̎�j�LOۖ�-!��*��CN��a�rE8P��8�/