BZh91AY&SY�js �߀Px����߰����P�{\q�1�b��	"��6���=	�`�h#�4#A��A�j��    � DB#F�䞍LCjdz&��@ �`LM&L�LM2100	"=F���<(�����H @I2��UbD���	?��]��UIiY�:�����Q�Y��k(堳W��������t�~��~���q�e�1s�
�;��F��N��?��$ej
����ΫW 67,!�*噺@�E�X�A)g�	T��Yx��]��3&L�"���8&��ٷ[$]Lkc^���@b:G8�����Ő3Y�G!����u��,b�$���ĠX�CD��R�W`�s%��2Q�0YՀ�4e	Ǝ�"�v�)����w5��H�����$�A'���4���������x�b���I�(�,�l��|JV�L�;��PuE[k���X:匌*��W�c��#���zc���_ji���̷�?��3���N�l)?tM��W�r�A��|WEV$�a�۫����sMj|�f.7�~�@Gb�h�ԫ�f�����|#��aْu��U��}��+H�QF��p�Z��0�_#�������Y���042�w�
b�2*��"�������p��k�����*��p�T97#���*�Ѥ��N�2I���8"��)���z�A")��ҖA�'��Y���K���z���w�L�	H�ALr+�I��4<���Җ�Btj��G��ʍ��8ʜ3��˞���ctd46�7��;t��p�KI�Ĭp��BM�A�t!et�&n�
��KI�����V*6�P�f!"$D���]����NJ��:c����J�*ZS&�mՑ�TH!q��ͬC�sL�p�X�y1_i��(���ߘv�Ő9h�jqD�Xyl���d`m7ݕ�H���M�[SgX�����BN�9Y���QX�&�X�Ơ�)'^:JUEG���5N����E�~��
���$͑�@��\��@��k�����,Q@����(�6[�C#��L2 ��U�g"-\���U�2*����w]�IY]�	���F���2d���O�]��BC@	��