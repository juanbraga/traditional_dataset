BZh91AY&SY��`R �_�Px����߰����P\��u�֤*P$�di�1M6�触��La�@Љ�T 0�0L �4Ȑ�� ��    h`LM&L�LM2100		O"j�Sf��� @ bh��0ԀUhD�  W!?��]���,H��\��)��F�{2Pb-��=6�X�$i`Z�>#���bt%q�]�	V�ċ���LD�I;��r#��p�j(@��AY
jiA�� ��2�[�T=����/�B	D�Fm1���I�!�i�й�KLp?�5��:�I�ꕿ��V6T骩K���3@�虴�M�(��)��G��lT ��E ����)��FHw#R�#yɦ��L���d���uJ�Z�5,�%)
��^�'P�7Xcs0��n�Ɇj�JzC0�GEko�3��p������ڢ`�0�Z��T���FA���Z)���yȅ���р���w������_  @ �4$8?�]d���:���fK�3T!f��Zb(p��r{P�� B�ad����j�W�3�bI�nH2��}���g��3_�m�O��g��������Ң��*t�lӮZ
#�&?�k�!7�N{	��F3���2�Q/2�`��#9�]�,W,ZΓ�MȟB�#́B��
�)���4fE�8Xn@P]e75�њ�vzA#Xw3�t��e�L�eas��VL"�lgmߊ��I��&�ꢋ��blJ
O�
�e��K@ĉq�9!R�0g,�L�/* ��2agE_�NA0�c�mJ���^0���i�`��y^cf�e3�Θp$+Ul�b��3�_�y��Bu�*'ۗAQ����b��eNVCs���7D�H���m-6'�p��sMP������!H$t񜡖�㇊Y@�2�p��V��`� yI�(Ba�lr�ً��Q(.�-	��ΨP����!B�9�IM�%�#��	�.3k��j�s�nD3�G	8cqh�i�S�%�p��Q�rꍣ���4�c��6K;I�8.�V�o�$F�T|bfq�̭N�.@��#��	�A�a�P�݉!�L�3Vvh0��q"�h3��� �Ey���"�v1��ಚ�2��E�<�'fyab,d���)Yi.�
eSɮ�E�C�B�:P=K�b�]�X����^�V9^�V	��w��xe�Q�ÒfL��\�Y�rE8P���`R