BZh91AY&SY�L� >߀Px����߰����P[pn�Өv�h%e=S�S�OFI��4� �d�A(Jzi2ji�4dhP  		4��5?�CM� ��h49�14L�2da0M4����$P�Ч���S�(h�Pz��FM�"��H�� �A@I�ˏ4��؃�d�?Rp��`ch��8�j����4�5�ڋH�>�1�����$�z�d��ve�+T5J�p�,~Ւa�ň��A�����Y$��Db$��	�����+�i��KnU������8K����z�H��g![l l�jw�U9YWgE�l��M႒��IW�3��N�̯U�Qhкr�ia�u���|Ͷ��'�,�)q��X�-I�(���b���4�y=T�H�Ʉ�l�8t��U��W��o���J��l�/4�Ϛ���m抛�}s?��M��_�>�k��}�G1$�3��p�^�CN���R!Ե���M.�sg:=E�l� �LM9��\��YL�5L���&����B&�N�~fuz����P��ұ�P��5�kჹ���$�<���r͈��y$vG2�d+W��kT��l0���q,f,!b6���h�B�L�aI=��)R1�p�
�u��
B�QZ��\��y0dɉ)��N������S"y/P�܅"7rw̆�Q%�aAx˞��.�NY�5��i�Vg8��R#�k^Y�h��e$�8�y�O�B[ �^�k`E���J�T�
"���T��	��E�JL�Sd�	���d*�7-)�E�%��B�[�Uq-Pd&	̤�Gt؆'�ϯl:�ʀ��O-�a�gh/ {L������K(�d�n,#��!&Ak�&G!�D��=EKE��J����S��Ts�z�ۨ��!
��Rd%j�k���%�\4���FS(EQ�(6IR��U�Bx�A]蓈�M����5�N����`%�&J�J�1;j��q���%@Ĩ���<?�ܑN$-S'ŀ