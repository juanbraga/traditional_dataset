BZh91AY&SY_�� (_�Px����߰����`?�� ��j�P��I&jS�6F���z=Pi��d���@h `  ��	�LC&!���i���� �(�  �4 �@  �A�ɓ&F�L�LDBe�����'��f��CA�M4<��I�� B�%H!J�$(�޼A���KJ��!��G��#IY����r��/}^c��=���)�o݉�=��?�*[�P`��wޚ����BU�!`�HT�X�Qԑ�YT�R:�;Q�֡-�d�|���o'ACi���p��	Ym�a]������� H-\�$�;�E<?g�}L2d͞0�Η!�nV�'����}���C�-ݐC�;A���w!w�Rb�2�2���I��[C|ͩ�zu�+ii��]�ƈت<]s���A�,��+��K 5�(�n����uEܚ3<���:�IZ:�3���Fڋ;;"��jTկ�܀hN�u!908�e�'Mb
�0��59��S#�{mv�4�K�L�w:��Q���nӼc��b�V1�Y{R�&��<�G<�T ״�%m�/VD3�A�5A�v��݆�=[�:�q�#F"M���wQ��g���C����Ӹ"]�&�@�b;��m�e��3�[����= �m��4u˰�HU�R)�NQ����zimUUZ�q$���
����L�T���S�E��b�gX�ٔ}v&l���4���ӈk�MA7�6��`� L8�i-��0�j������f��e�$�#'�f�G�A��'���5��y����0��W�&�����X��B�Lb�@�vj�v�dЁT�>���vF�#JNi�wm�0&yz�*$��(V^��l'y�}!l� _�ل뿠Y�����ar"�2ZHEY�w�ӥx��ô/r�k=���l�]9�m`P���WV�!�l0��O��[	o�a=ʘsA�G-ʧ�c�� .q��(�B0��;�N(��Ki|qz�h
��*����S%My\H(U �1��X{��G%�xq�@�S�)��P�h�ӡ��Sa��u�(<��r���Ѭ��m�q�N���i�#m1�{�˔��לнm��k0$���p:�J2��.:��@�<֤XZ�T�aENP� y���R�$(S��f^�!D��͒�&w=@�3W+7-)�E6x2��(�:"#m�1@���4^ �s��e���D�7R쪰2�U����Ӗ��u.F58�{�1]F0@��:G�p�9�����u
��KK��Jh�%�$�0��c഍�TZg^�]^*��V�����e��gpYT�c� V`�<[���n7#sP�ir݉~,����e	��4k@232D֮�\�Z��f»Պ�FsvwhBkt:�jR�ㅧ+�ɀ�o��7�]��B@~��