BZh91AY&SYSrO �_�Px����߰����Pp˅P�sl�����ICF���
zCF���4hh�jz��Pѐ� ��  S$Қڧ��OMMHh ��@���a2dɑ��4�# C �)�MS���&���MF���i�� =M C�"���(Ȣ\�,~����G\.(@ވL;��D�T*�V�J,�t`��|�s���I��n��Iq r@��	����tp��Y/e�B9-9�1�s*MhU��T�E1��K&��P�^��#ĝHe��tXu'����'4��Vs�"f�<@&��I�g��?id �&k��x7��rk��Kr8<��P��k-v�4�p�LdWG�;#�6A���B\�s2YY�R�"HQ�q H�A�E�+R8�H!���V�2IDZ.A$$�2[�0�w��
l:C�%����D}� ESӵ=�Z�uhP�XaJ�˟{��~�{|�d���X&���O^�mM��b�}�[��*֒em�Hi2 >}�^2���өuO�wsg��E����3�	-(��n�� DR��)0R�F��C,;:�[/5AH�zw\�5Nj�BD����D�G?:���Fd��G�G`��62������M�q2�3�T�Z[<�?|^Q�$�A'�I�" �ON�8���Py�r�<��tYrܙ�u"0��	%v�G��A�\E��E��g`�&�P&�32(�Q\�L�@dcs���;����U[�F�:�3���w$w��o���}q�E˅xx�uF��8glۏ�om����Y߇��Ĭ���ഇvYq=G���U��D����h�g3�%-�flo�!C��.W��J?��5�"�U332L����� 叹�G�a��Fq0-�t� 03�i�vok��H��P���׺<��{T�l�bC&&��禤�B�SA���f�j�pn��i�/;%jVX�ä-
�N�T�O�s�+
'��1@AR?z׈t���>��͏B
�釭i�jvO��Xc<
�n�:�_� �I'q��udXק�vHH���b��'��g��P�<�v����A�\D@F�@����%p1�v��0"�A��G������Ge� �1.���R�mЉ���@i1Y���C	��9KUR�%��ͳ����g�De��Sa�)��"������ò�r��U��`�V�l5��@�PB G���dK�g49�	D'�:g37Τ�s��A�U!��%��C�Lv�N��]տ�:���$� l�:q�����S (*�0�,,E�1"�gLb��j�a�樊&)j$��~U�0���V�9�k;�a��f\��^��Vi`6�`5fVy[,�ܑN$܄S�