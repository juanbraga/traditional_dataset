BZh91AY&SY���- {_�Py����߰����`<�<+�    �    ���Jy���M@      S�h
��� @    �R4�i���&L b@T�Q�=A11jh�M!�d2dɈ��	�����$@A �2i�#5&&&���)�8�bH�d��!,h=�@������?��Q'� *Z��?�*�����6JD�T�I�0Ėa0��0�d���|sOBx1�Y��1���i"�""""D�����(Z�"�Di��"`�e6�� �m�B�!B�m�@�ؠ" !�n!B(��r�˗-h�l.�ɔy C�|d yc�|�#�;��^�A������!�R>)���M%^,��R�os-�N�r��wQB�Ő�t�GR�mj��#kR���
FCX�)�T	���WSx��3��a;c]�w*舂�j�,�P%�m.UZ��!R�(�%aW)k���x���\-�\�Fm�ܲ��%-���[y���S����G�M�
�B@��k�$�c6=���aB�nY[���.ޱV,����Ɋ�f�%�$D���DDDEV�Y*�$DJ���l���h�Ubɤٳ����ۛ6zᖾ��r�T�QR��~����V��µaft)��-B�����ə��$pN���<�@��$R�MZ�M1y��b"""""x"R����&����?T	X͵������������.*�)���9�YbE��nو̼����x_�y��o�mW�>�g�������m��}���^z�W�G�Jڼ�Xg�D�ƙ�i>JQ��'�r��λ�0�m�9;l+r(��@Z�ʊ�x"�v8׿ ]W�y���7o|�C&6�m��m�������u��F�i9W��CK�j	H#��T���T%p�(�lOn���I���p�ۺ�rE0:]MV�$Ld�S� x�f�tBՓD1׎�m��m��+̿P1�>��Q�R2 y����� J���ܘz#,�Xz���J�,�ܡ�o|r܋�	��d1sw:@�/��5׀3>�uz1ہ,�}��m��}������z��K��D;�>��s�MH�׽��F��h���Y)�dWpc��R'o�@��cp�LSL��}��a�©��Ͷ�m���E%�S�2 +6!̕�OS!�rg�bg(#��-뱣�7�W&�R�ɉ&g7���f���7�����=���r�ƈv�[ �#�fT5��m��m�Δ"F"9R���x�0����C!�u��Y���/���7y��XT�B5�-����̈��W(eozF��.<�P��3In�w�6�m��b:K�w4#�J"x�Mm�eژ���w�r������-R���0�[2#�t!���r�R)���m�(����-��m���>�R�r�A�h{���q�N�Z�B��q�krJ�<q&
۹wRͯE�U��ZS|����T:�4�{�n������\T���3&8]�S��p�m��|��^�о�v��u,s-��"G��:ʋɉ��C���1�(g��;-�X|A������;S�w�JU)U�UR�� Yf�s�.�^p�=�wefJ�W�%�н��R��T��X�QJ)W�Z(�(���R�QE�����QJ*QR�QJ(��TQR�H���T���5��E��R��.�U�?E�d��RL.XKк�`I�U7.���ʦ2RՋb�Ԙ�ʦ/Y��,�U$
��*�U�r����uk���z����}��b�nY��oW�����L��u�:�zp��?�K���]�"m,��I�|=�i��3�����\5f�ze���1�o���sS�vS���szdɪ)B�ZR���xH�m����ΎIĻ�,�d�ZL���1p�%<I� >����j�����Ȧ�x�]&.W�ƅ,��S(�{��뽬wҤ��Kli���y��?,g��0^�Tu���^����PeD"��V�W�tX�4��-��c�}ċJ*PJ�R�B��I�7Ri&o�o�&��н�c�nj��̤��-�@��\�����������)b���,]��Z�y"���x��4r�7K}MK'��2�z�;[NwS��1��z��lߏG��!��(�&�%�v���2Yoj���t��M��t�����(xټ��a&�8�82���������V��')�,��ə��;�ل|�H�0�i�:h`R�O�bݬ�dy��̪�Œ�)i��k^�Ma���
LaZ���i+�����H�]�Gk��9��c����>~�Og4��F����uʡ�E���z��#9��$9�0�.����' �Y$��IR �yqf�7���wc��q�{(ӎ1T�Z7IJ��tLX�+|�gR���#E6���/&۵�bi15�d�����Sfʹ� 4T��[�qM���Z�[{�[��V��r*-'�$�1�6���C6�x/�˱���C�1'��%G����ϫ�h昜֍ӫ����7�O[�c�铝��T��TQ:���{?���)��?9h