BZh91AY&SY6U$ G߀Px����߰����Pѡͻ����&���I��MOԏB�4 ���<&A2��I�C�4����#F�h H���M4��ѵM h i� � �`�2��J(��        $W��U� �E��I�����c�A�Q�OGV+A݀�� qET-(�mPTx��w��]�+ �~ȅ]�4:�2�F[^>��df{l��1�
렑ޱ'����U��!+��`�k�]�ѯ�<7m4�S�v�&9��,�k�>5��N���\1�o�JO���!�2GV�e�$C"�"�lv&�W)�K �i8ڪ�h���
�	P����z���|�llm�����ҧ�"���b����qh�f�lab��*���	��e�P�؂)��>c�L`�t_w3�S�Y*׏<�ͳ���^P��#�������}�.*v֞/�����]0��P��=�����NH4�@�aTOs�C�i�����8�ҍw!���҅��+LN7]<f��*��f��2y"b}�"|Ð���$HJ8$��dd|m��L鲛n�'[}`�A�|�szqY�/٥���@E_&x���wH��MR�0�;	�%Hq�	ѳ��=���r�_�d8�*N�XJS��c��F�#jpbI���X(M��)y4,�d[�	����G��ʋM����Jq[�e��^j%"�I!Y(h;{��8�x�Z��з�fG(��h��fR����b��,䢔T�Dh��$��N�P%&R�"N=���R�-�G%AyKf�Lt�R��3�mk*�sy_��P�]�9S?�;0�)�GC��ו�0mP��\@�m<�%<cH�Gn�-ɉ��@�x��e)��f�Ldbn��)EX��5h�R��C�=ZM��v���o�� ��X^V
8�3�:�	�K�P$Z��>x1zg
��M[�Z�]�a6l���Ĝ��;H�`��O)=
���Y�C�V����Σ6x�[I��7�d�_+���"�(H*� 