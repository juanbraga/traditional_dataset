BZh91AY&SY#=�k 4߀px����߰����P��d9�嶖�g	$��H�j=��z�M � ш5OTz`�z�C       ��	2O)�#�h�F�A�  ���b�LFCC �#	&���{J{I��d���@ h����"H3�'�=˫��,Vhѐ�i����,C �GCP�Q���>ď��Tc��tlׯ�P�b�h*� �p�����5;�%I�y��+�F�C�3P�W0�:I$*�T�E���iѹo��m4�y���[�k��{cB�.i6L��!q���u4�����ϴ
�Lq�7�B�e��� ۂ�A���9E�Qn.������~f�`�O5���:��X���M�G�e3�L�Y����)�����Y�������Z�U�7�1�,��gJ0��k����Tl}��������y>�=���&�z�G�����X)��]�+�?���z�a��y�&)���Y�o#X��e���d���
2�[_��mJd�	.8-#�^Z�)��v�7���FPZ 	�\+AQ_E���> ���O�lч%�F�=*�E}�1��et�PN�j�Ƀ:�s�6�gՉ���U)�:�1����b��W�w�
�5���zP�ߪy�zr��X/�+�-�HI�l'#D�"8'���5P7|EM���jG�{�r�լa��1̹i>ת���U��]q�hX����-e���j�x�A�k!�A(������&��15��T	I�P;�&s�ߪ�J�8�t�%5�j������g���9��9Jū)2 ��b�5�b@Ɇ�)��I�6����� ��r��%\�Ǣ͢\��p��m�!e�����=��d����tU��G��&�s˾ve���H8��T!�ly�$ï�۹�a�Ȍl���"�;��2�e��aZn�����-^FE�b�˹-W,!�<!z)%f]e
�=�J�L��k�o�w$S�	3޶�