BZh91AY&SYb�* <߀Px����߰����P@{Uݹۜ�XIi�FSi��T�z��� ш=M �@�jy&��h��     ����B0M�5h� @i����&L�20�&�db``E'���4��LCCM��hL� H�8@�$A ��@������T�+1���ê������5��Z5;cq4ƮX��v?#��a�m4��+t�?���8�F㽒T�c�}�H���|��6��G��	V��$#�xrX��?Z�m4ޭ�ȳڪz�ϋ�7����#����7N���*f��y�����X�`�)RX3�J���I]T��^�C�2Ӎ�{5�6��ߙ��4�d���)㔼z�X�Z�fQ�l�bvf�����t��3�;Pd:�0�Vj���D�K �dz�^�Z5��mQַ�{Z{�3���/\�
L3p(���Qr����;�Ϥ��>7�F�g6͆}�1�IB�lEr�תf2�[���cP�0�q�U��z4�)C��!M��K׀�&ؗ�Gx~��Ǝ{��d���#�Z�dN�t�Qh��B���(�6չ��6���(����1�f�R�"B�j�Ɇ�,'r�E4�fy���𔎹RQb_�B����4��LG�s^��$����bїt��-صHs��ѕ$�7밼�k Ej���1SZ�f�G�d&^����(�E[��ď����2)6������q�wK �&��!t�#��}7B���&�*%k�Ap�)V�N:`#��3:���KJd�A6�j�A"D0ѿ`���Z͝$�³yZQ�I��@�e64�VQZqf��L��[ c��h�;
h��Y��K�2\,�Sl2�!Mb��6��xw�)FW,(T��T�ǻNr2"��{a])ئ�jH�9�Q2�+�@�v��
�
�U.F]B�QQ�%&A)(�,���'���P�rP�c� V��ފp(�R�th.��ݨ��yKT�NvksSA����ݼ?��H�
]p�@