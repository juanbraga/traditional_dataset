BZh91AY&SY��{� _�py����߰����`�x>s���a���[�`H��5����#L������� � h5=4�2��  � �  *oCJhS�   hi�  S�B����� 46�h  � E�����=54dh�j=@�$h�S�5L�$m�#F�   ��!5��#@	Ht����R������`[H�Tֈ�K	�~,�G�3��,
Y�#	��t7޿�;ցT@TA�XQ9��2HN��4Q��'k�Ywe��5ʳJ�El�q�Η��[Z�y�Ԡ�j�t��F�M�lLMQUSj��4O��0ȥ
Al�T�/�A_��k<��Ǝ-X�a��IHۚ(	f|(���xc��b`��!6�@!�6Kw��SK!fI�6g�r�Sf��������d���ͽ�~�G1�����˦mO}n|a�.(��>0��Nj�+rKU�qp$�lxH�8 0�v��%�6m@8��}Z]˰����N�t��o �0� �.2����&��� 別���q[�@ښ����b��v��ĶېZ�ÓN-QDN�wy����:.�$J=Z�]�)]��TIfI�U��ӹrp���+���*2��:3�%9T�Ӱ�$�ɫ�U ��ɎD���@�j��-K����)r�M��MI��53gW��
�Bdj�K�b���L�\���i���et�w�k֯SF�snm�.'�!���}Ɩ�,Ͷ��������HT֭Ȫ�6�ސW�Γ{�rw��8���+�� dKq�vb+�)���(�3d�8fl"A�9��TԤ��$�µ%%	�c$�+�ɄS BB�@ETG��2�9ɂvPdO�e�p	Y�����;���SEUoa��.Ķ�%��Y���}����"%T�X.EM�v�y���ƻȝ�V�L�80��@��8�8�
{�@|��mN���GaWt����!:VT������w�3�*�гF������X@i@����DNGa ��8 nL�W3ǉK"	���\���ۥ8��`�o���݅.�ߑ�Ǌ�c6D��nmF���$  �3��Gub��qоG������/.,zR%���{��t	Cw�rqt5�Ϩ.[�<�]` �q`*"%��H
:�k����]c�?ir�P�����u�\��v���������5�p�d��,�/B���#E�ɳ��uJ�<����7���@��ITw��6�a#���ll�hu����I��8�k�q�$i(�n--ؗ��X���|�c�y���P�nm���0R�!Kf�6�R�D��E����b��-��r���Zl9���<����:k���+"���s�|����g%�ZA�{��PְY�f�2�D����Yq˵�ri�r�)ܵ{`���dӆ�ʴ�V0903�X��T�y�V<J�eDfM=t&W�(S���BA�,����:�c'��AY�Lb�_|j�a�5�C#�`V���>��b[��:JmEJ��0�qׄ���.D���Q��jd��V��U�ܑN$4w�@