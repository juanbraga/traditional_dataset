BZh91AY&SY�\@ K._�py���������`3���@r  � w��M{a���z�(P٨��-f5KM 	*�j���h���ZF�JlQkI w�    ��@*I0� 4� �   "����i�&  i�� C��db0�`!�M0�!�F��jy�H��  h  �   i""�F��Ѡ i��  I� B`�zS2i=0�z�S�AN}�.T�E�ߴT4��T� b?���*� �*K�������1�BB2
��EB4��^���.�*Et"�FD}��-C����r���=_7݆����EI$d����VIRJ�)"�,%d��VH��@R P�J�+*Aa* �E$RJ��*(��d� �a �H��,"�)���XE!*IPR�,%B(��RAm�# ��Y$�P��Y�EdFA��%-A����/���<�	���>)�G�;��1����w��c21�MU*�8��\1 ���s0eF&��BacV�9!\H;Y0�S�ۣV��Iպ�?�8��������۹v���D:)L�pjl۶*���s.g!�"P9Pn���p�#��,�BbdL)*m�as'��偙p���%�8���P2�&�f\�
 թ�*��54qK��	]��a$��2�R1e)���JTNE�y���
���P6��td�x*n@�Xg,J�SB$ui��Vݫ��p���L��&j�ͩ&j�Ybļ�4.�J%5
x B�3"ȉ�3�b�1�ZB�P��f��(UC0g�U��l��(X� ͼ�`V�[�"�fU$�rSR/�1]���Z��)��*��Ȭ��n�@8���QEK��J�෎��w�nd&�(/*o�X�QDeӛ�3�/$��0��/��̺W��Ua/2�W]�� Z�qR�70qȁ�l.*S��91-\��!Z�cT�T�w��W0��Ę,����� �b�U�T1�_�[���^��-b�ws��$��d6���""HG]Y���Y]7WVn`�d��o��ןA�8�p�,_h10/�y	_(Q�i�Sr1�ٜ\K���ՉY��н�/bK^�Ne��Y�t6b�൳G<�&k�-�@4�J��LMf�+f�6�[.ZJhKp�m��(SZF�׈�q!x�(���,�&v�R�HF[5/��Rk��.&���
�nT�[]Ń��|q7R���RjĐ�i�\�ĭ�ګGR��:�-]u4�]v��&]�h�T6��M��f9�mwY�tb��fn�oӛ]��\����5��A5Q��Z��)"��l��]�ƥҍ�`�T	��I�5�̘� �i�V3M,���贱-�����i�i��3s	��k�"�h&�atH!��vm�����v�X��][n��3K�i���ƭk]֕f�q�)kl(�7N��^�v��s+�T�m/,\Zk�-\��6��Mf�`M��k�Z�z�8X�a}W�"��2�e����/`2w�=�jT=��D���2쇱��<fy[��[+U,�8�
�[�ʼ��ECT[N-E�,N-xB��v� �(���TwLݮ���iX
��Շ*UA�Y��)++1���H��7�M۴Y*�aq"�aY�U��aSi���
�)�5�BlAL`,PQ�*[u��f�I�aX,PU4�������[j��G�M2b��E�(�J �H/,��[*b���B�#m��,��r�+:j�0P:&0���R.���\k:l�f17���1�YZMu�T7�����ꙫ�T��YPK��a�
��]���1��*j�Vsv��:8��Xd��6���m�ŗ}n��R�P��G�� �� �FJ�}Ǯ�A�>0���m��kT�'��s@æ�c��tZ�%�J^+n������NRMC��6����1�WM	�&F!,�å��64�ldج��.I�F�X�K1
P���5�9Ƶ�6s�F�Y��-��M��K�ܐ�8H@�A2o��8�|�kWY�aR܁s��%,�WT��ޛ�O7R̤W�tDeUystƦ�[;��r6t�Gf�}X�F;7�^K6���#��Үz�pj�r�2�h)�#��r���:S2�9�s*��Æ�0�2�[w�q"lg|��4��)���023��	��V`�94+j4�i�tlPm�]4���â@�h3 ��B��Sl�"t!Z�m�ȍۺ���\�j�S���.�cȕ&�����D��Լ}-�-�O�v�}�[XƜ�F����#,�pjUD&�8�֜܃/�Ϊ��=#d)	�;nIݬ�W�ZV$�.������@�y�n[�Y�sL��02���F����']=�V�yZP��r� �E�*�Aq7;����:Dڱq.�0KZM50�$�p�l0�;�.���9"�	75Y3�jq�
¾�y�!�|j�Xc:ofF�^�e�]m�ALMR��'3�ИjcFkv_j�2s�oO�
���F�*����R �KyS��gț�sEln�uJ���̙�h�e�;��Yp���_[UP��) 3]�
�iX��Il���>y��[�h�������$�i�ݼ�mo�����{ݒx�f�b�N�f(Emc6kң���S,_�WƎ����v�^���k�#��J�fYӾ��Y��vV}���U���Ad@��m��c�h/��['M/]�i��z�l���5���%�G�n��L�]���"o̸�7��`eJ�4��戫ڤr�P7�*E��]<�]Z���R���0F&�ni:.pѾx�8&fl�˕��wK��+�&bRaO�DkK�b1��W�٪ƍ%��q!9@�[d���#l�T�Ccg�锂�`�
��-���g$�A��{���ˡ��L)J�@����� YF8�#,��T�)S\�Oo���ۣ'}ȍ��c<�@��w����>�j	�T��)�Q�6��Rc�Z�bi�S�3��C\�
t�-"��V�v�z&�i|q��&[
��4ׄιBR��×�cU�
Y�+�^�9P��\/]H`Kl9Wft6���yc����Æ�Z��(�u+<'F����-��V�>�4˜�>E�cp�`�P��R��2��B�� `���~��4��Lx! a5�=I_�a$��桘��p7`�W��^�θ��d�lI��s�-{�F�*Z���6$���H-;�/n����bCr� ]m%HE)���i`r��X��AJ�3lٱm�ʱY�7Km�6L��,��Qe�f�t����hй�_Z��ky�=[�I')&�;�ɲ�9ք�.t�Ue�R\���t�zJkwpݮ�@�-g�5��U�uڼeV��1J*RH���T<���!9�����g)�Ì5�/��,���&r�����嬂�d�.v���Dbqa�;���a	Y�����V�n��fG����/��@j�T���]�����K�S�Ǚ�_S����b<a��o�[���!P�u����psf�Jg�c]�쒊$)�.�Z���|�.@�a�e ��`�b��A5]��\\���Pmh��j�F�#k���W���o�R��0އ�Ay��P0�p��c����&�O;Iq��a.�Z\o?(~y7����3vb�����E/2�/N���~�f2r�wʼR�vFXv��2�"T�m���v���ːm"�o����e�Q�����`o��렳*�T`���ft�P�߁�Ŗ�Wm2*T��3YoPY�2�
���UL�����&2ҡ=�|���o[�f$q�c%�V�A	 Y1���-I��:FgS��S�rf Ss�4�S���f�OS���U�2c�T�,�����eTs�XX�$'��eİ�w�gV�&�"�m�	�0���;[R ���#���u�U��-��۸̍�Ȼ��Q��[x�3Sp�̭��]Sb����nuX��]G��<��m��c3;K�i^z~�X~�%8]���o��|��S���![R�yM�*�_��M��f�;}���!
�0���e�� :��M�L׳2��&C\ ����Lٯݤ5�ճ��;z�z�oixVb;	�f�0��tdc��aU�q����W�w$�P�J'��*��������&/���2ȼ�ySɎW��@쀎�`�����>��jZ���!ޤ=�Y���n0v�JH�xFvt�������2���ɖk''��ӱl���82Q/1G�}K�k��w��;ivک�냫�^��4�"�j��p.B��jN��TM�ͷ�����r���������Θ�
kP�,4���^^X�ɉeH�|uіu籏��a��{$6�q��FZ��8��S�mi5���m���+<�ϓ��	fQ��,��#_�/�hT��� ��`{k�5�Y&s��Ǯ��$Vfzv2��\�L!\�i��BӋR�MCEm�B8xנ#K��O%�y�����UV��>y����"�!�,���_$kv�G�hT�����
ۭ=ӭ㯕4	b�ɚ���Ҟ'gϝ<�������ƾ���2T�-���=�� �{=��E�D }E�{
̊�[wviP�V�I�A	��ObB3jb�Qr�ԂȺ��:S[M6A A�θѻXf�xf.�+Z����뒵���(�g��]7��)l�GK����[v��:KqL.Z�h鮛5f�auΛ�T��9�{K�HΣ�^���m��	f�
�dC8�]�6���*j\��:<9~W)�Q���%p5$�y�S;k�sB��(��7�l�k�9}q�y���y?�NM`���N��
��Un�6:g��M��\ ��y��d��95�������3�gB���;�N�R��n�BdWF�B��WH�n��u��8U�=��cZ�eN+�}^��<����Q:�̚=.���dr�D�6�#����˓�Z m!1L����M��a�\Ar!��Lĥsc!5�A��^��k{���6mGn#]jY�6D$� �kq�~ɧ`�V�L�%ظ�:�)�ץ��lW���� n/��~��R��b��n�U��J��uIY		�w)�L�㒮��h�]Ӕ�$;3\3��"���hh����U����㵵85H�<dt@��:f�o=�Gp��A�Co{=����Zu����W
�HF��r-υ�U���YF+j_��47K�މ]�r_�g��.�j1{.�%�l4����0E���f��<�S�{�M��@�dR�zm��F�l�H���`���"H&���e+£���,	��tߚMG0$�l�z1�^��>�X���s,�S識z�3���w`��o{��^�0�;�骪/��Oo�{S��u&����"�FXZ?3z!�͊��H�"�Ҋ���iT�&j\m�U`��	ϥe��*�\j͚�p��s�;L��3^L݅f���f.&��.��^���!�j8V��>��6l�ܵ%X'���̻��Z��C���ٮy� �zvP�o/�r
�W1�Fl� c�&��Y��E��L�Jkt43-Sjz�/K��ן"&��8|�Reۯ��К�a#�� ®�!3k,��nǎ�S>��0]�����q��D'3����L��-*A756��D!Zjқe2o;F�7��.6T㥕Q���"�b�Dh�F�rȱC�ђ��%^�[}=���eM �f�q�ҏ^F��Mh!��j�pvl����ٙqWv�P��PJ�*�"|l;�2T)s7�fi�� ����J@#�;]i���c\����;y#�v�Ȝd<[�,*�9+.^l�LM�JK"N���ۨA���!\��F7ڢ��m�f�w=lP�.�����&F[>��8o�K�� ë��sZ��b���`���;�Y�;�����+szn�,�x����,b�}�L9�>t��^��e��f2�9>z4G�p>�-1�d�4��{.p��I���mg(�a�P�yR�ϥn�8M4
ܚ5p�"v���`ʺ�;x.��!��ta)�-�fq�u�_[3�X�RW��"L�c�P��DĖZA0�M�ڮ�L\�qb���23<]��\lb�:�d�f"ʶb�55MkǙ�1��3V�(�q]�`�w�N��N����@u��rd�8I&�E	���r|�J8?{�^�;����/(�I�rn#f���t�
fÓ�A�M=H����p(�Ok8{(F�D���E�!,̘����𓽦�u33{XV�O�l_������E$I�~N&��S(�o��t�a�5���5Zƌ5Sk�i���$f�����I��x:m�������S�����:��.���������fr�SF�WjI�O�B)�TZ3"���\x-�kdĹ�ռۀ��&f�Y67{CQ�S��.���YW��$���}z�z�_� #���{�+���f�Nʼ�n��A�2�8O�Q��՜��u�dzL����5U!�FT� O����( �����T�ްb�-�=�����kw! &i"4&D�pY�f��4S2��*�L���ǭ�yi�+��ĤO5�i�nڅ/�I�&E��/�w�y�]i�oʟI��x}�bz�F�����P��cF���N7-�1���ul1�BT��'C�$чn`�H��N�C��XÁ��59�Gr�*3Xd!�`VK-D�3UqG�G�}j��ö�kf�Z��Tg��w�ΫL�G����p�/ ������Ig.�>�GG�A�����S�ݗ㖲	�`���=%B:�[u1Q1[��&�-�	�.}�`�+�q�����s���q|�Yڞbn	l�f]�Oe`XVg�_�<�,�*v6hD�ce�����%�4��=�g� ׄL��n���{˝I>�P7
~�\�$�$%&�� �� o?
�W�B��t�`%�4�]�/�٢�=�9��x׹ʊn��=z�w�ޑL�]J�m����JN	]���!-T�+%79D�'���b�:S:���g����auԁ+'�Bf����b���VN�0U�Y���V5�C��try�k����.	s�3AhO�v�BID�EN�\������+/��Ĉ���1t���KZ������Ag��Wb`���U$��z_�ݨ�T��3@:�J��BڡT�}��G���1��{�UBN���jN����P���T��?d8B�  �  n	���i��(��!nIc��G��lۜd-�])��a��t��5�l�\��%-�]`�+[\ThE�,�e�/���'~����wġ��k3���-H�S�������҈�ݚ:�@��sr����h4��p��E�S��P���Tg���������ǥ�"�����`��w'�-������E�>#P�̯:�4��h)�����׵s���ܩ[� �j����X$�v�1�l8;OևMi�Y��U>9!ݤ�佯�^��c��4A��"���	�H�d�C9��b�
8�I�h^P�ǥWFzc���^Ğ����w�$ߪ�M��Uͮ��$!k���5S��v}�˼{�kf2��g�sl��+|���3������b%鱞�v�{^�x��(t�N�gim��KP�m;�1�;g6#:��{������`�������}u�6�mv�ղ��T�p�6Z
#D��J����o��L�9D54'1����̙�NMYx�n0Q�ΟlMdH&�%q�6�/����5v�i�8��r-DA1�g��˛>d����^	ْE�-ѡW_@KQ��Q�*����o�x:ƽ蹱���̑%��3��1�C�S5���j�����bXa9�Y�UiQ�FOc����g\�������ϯ<����Z�� �^f�̦˩V�n�W�%}���SՏ;�e��̧n�ZH���|�=5�vgf N@}���7�����fA:��)>T�C��ާ�^j�O�
NZ]4M���W0@̊�Z@wwۛ������l��;�,�Ò�~/sz�Tܙ���@0 q#>����e|�Q�$���ѐ��٘�cM�1�	i���2`6K 4��~����|9?���n�H���v�y`�3ﶋ�e	�A�!��E�c�sۃj�n���ҭ;e9law^j��W��nnn�s!�vex0"<sq�a�Xه�r��L��I̾�0���$���9��@�%~7h4]9P�uﺥ�,�Om�x~G��|_P��H�/iU@h�$�������-�>��f���1�"����Q��z��+�A�!�D� � �*�T R�iR�ղ��&e�R�
���%f��H�A`@
�*I�4b�`�6���\$:��Ym��#*L�c�=��H�\�&��W��|X����n�?�M+���6��������C󍿌l�L���bn3?�oϯ�����z]��<;�>_��r�x��]�~�O3������l%������[��37�J,
*�������O~E)�N���2�~�6�! EC�H�����u�O=�c��/$��z���.�[���~=Os���;E=�?��g྘wN��0����
aпM�v� -�/�NF`?(p�c�2��(i���Yn�N<us�����T-�{��rȻ��1��r`  Ȁ�%�R@DP-H�B"�(��B�50D��0T�K�~�e��e��]��ñ��LsC��j5�#FIg[����/2��G�Y���V�E{����Lbz5.I��0~����;Xs�s���"���C��g�M�N������Q����m��i�j����A��o�0;'߬������ϧ���W�T6���9��J�����[��}��鞏����  ��P���~�x�sϛ%�'}U��]4f��j�j(��,�:�TA\^���Si+qtѣP\�UU
)M�`ya����1KM0���)+�`fN*���M4Mp"br�H�&G[���!:��rN`P��1��N_��M~8���~����<�}��&��U:�>�iP>w���'��}��ȴ �N�<|����z���EB����.}Ϸ�iӼ�8�waÀQ�=:��0!]���L��KK�i���N�;�g܆�:�̶떧�����a�.����1`k�0�Gp�lNv�sy�7����N����46.�G�n�n�Vtۡ����$O�ݴ�E���M� ۇ >�]um���M�J!�pK�Vz��0�0�2����2�?�.V���@�1�c��:���)�"� �