BZh91AY&SY���� �߀py����߰����`�x9ܰ  ��UE�$Dɪ��=M6�������H� 4�����~M*eOO@ �@  2d�L&F@��M#4i���hS�4�h��i�4�h =@8ɓM0�14`� Ѧ HMdjb��S`�� �� =Lq���l �H(^�XH��y0?� � �3X|�	"�6d.���۝�[�m�v:�,����X�4�4�%�%��4��T,,���I��G��(�vE���x�=�Ke��������0|�gˤz�dK��p�Phd�Ęb8JII���pũ�L�Z�V=M�_�v���޹��{������"5疬�*iӪ�
dR-�� ��)���揜���I�j[�;1��}�B 6�sW�G�NC���7�3�%_C�lj�z��H�B�n�g�"*�bcI�k�cL����OCD_4���x��(���<h��w����C;*#l����d0M�EZz[����昺z.��A�>jl��gJ��S+]��5f�6e�#1p��>#��
�Z�,�eW�����o"�/&�QQp�wRgo��$�S�\T�S�M�����������%��;;xG�PN��Ǖպ���ֺvy����tM]�R�L�D4,o\S��v�L��I��Fpyt� ��Б
(Na&$�K���3����(b\:�xeuO�Q�r�ϯN�n�!�[ą)�g�{l�*��K���6��@��&ͦԻJ7p�Y���պ0��Mmj F4�U�A��Y�� �
[���b���и�K�5��^@��G���L�ȷc��w�3�[��at��*4���mB4(k*�Qx���N�3q-	�y�l�ٴܹry�d^��\�5<����\��
Rrd6:;S'!4\���5,��q˰|�QO��"�ݤ�M{*�C�e��_�N3����l@�Ç��KpY�O`��x*�K>*�o��R�kd�H��B��J9h�D��%̍�%!k%$��!�a ���^F��Y��2e�v���@6�*l޽|��r�3�M8����{d��j���`>�U��zi/��r�]V���wWEٰ���Z2�tFB�ӛ���3/Ð �Ht��K�6�d�a�ĥD4"��!'��GV���6�Fşx�mt�D[����U*�v�c�o	y��i1lڞV�C�����g?*�#}��V��O]��������`�o�Xl��&-�(�V] E	4�f��<<���4�=B@ +�^@�Y�K�J��n&��T(`�S�9�W��^-�:�$8M,8Y��:���p��V�d��x�h�7^�E��Gg0�;�e��cfܬ�;� �������̩)xN�7w2\N��A�D��;@�K��֝��2cqQ��4�4(�#~���I�<F��D$;'�Yp�eF9)h�OmJ�^C@�L�+W1��Fe�
[)�i�6(�$�1qË�����ű
$Ϩ���E�L:j�7hniv��7�#o�!n�Rc���i��)"7s�0N$;��s�7�	<)Y���>]�S���ec�W!�U��ȥ��c���R���ĝ��T��E��FQ��h)����3fݔ�6&D�MD���Lu[uãnۯ�ׁzB=	E24kHx����߼�7�8�������2�{M�����tS�G��?�w$S�	H\^