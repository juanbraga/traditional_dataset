BZh91AY&SY{BE� <_�Px����߰����Pr��鑶��IIFG���?$����&22��Q	��52��� �     	Mښj�I��L�4c(�F�4����& �4d40	�10� ��ji=&č�z�2m#@F�I�D�y�
1"B\
��滎��	4���!���7�0W��ml��AV�\�&}����!����ڿ^��yE|����D�G�Wh(E�o�v� VsP�Pɯ��nV��IH^�x�Ƹ.��u��ci��w�Y��ݲ5�:�"[�[l��h�a���@̕�AC�ic0e��Y0�Q`��MoD���Q��{�攐���I$	����M�_ĔL���$�F��2�G���!u�(7��P�Y�AD���/tpʍh�G����f���ot���f����o�:�LK�L�ɝT3��w���]���ۑ�y9�6B/����.�D���
�;���m���8����aa9o?\����;��!�$�S���� ��Wr��%��tx����g1�l�-�{���(��ʷ��c�8�aF{V����M�l�1���)7�P��P�H�9�S���A�s�O5�`u�/Wh
����Pc+�݆e[E��ה�\��9V�!�������`=0�zi%�Z�+�h��w'r7�J#lq=R%�n i��N���\�c+m1����?�U��R���%���v8�k8�@�BZJ���0�{zB*͒�P�ZjyBh��%j�(%k���	 d�!�vN���>�0T1k�'�0ȋ�ȗ��b@NR�m�Cqzs"Zz�E~si�):�7��c_�
~��s"jYZk8M��b�la���-I�������t����W���%IQ
�T��}�P5��ό������ƃ!{�Y-Sy��0Ң3WQd�bFb�D(�����JJ7]��m�DDP�r�+K{��F��ኜ��z(.��mʆe�,P��c[ �ɐ_?�3�ܑN$Бt�