BZh91AY&SY�1� �߀py����߰����`��| p  ;  
  π         �׀D     z @�/gGUV��-ݠRE� �M;a�Uu�Wp����GmUG]ګ�&��P�@S   �h�l 
�UA���*4�MPI�����H
  �[
��6�D�f��t�A���`
V����m�� �B� 4�3U@��� ���� 1TV�D� @S �M��V��0d �,`j��. <)V @�APO�T�C@a     "��M	*��`      �LsL��Lф�hшd�� B'�RM
*4����  L�4"�4L#2i�CA�Q���i!)�D����1����!��5g�S�"|'9U-V�b"
�_�8�D��TE$��
���I2H4��"��'��i:dH��	"���a�e�C�z!M�'�T� �����N0;g������7�5�?.�ۿ��b �a	"�P��
I`� T,��@��I(B,$PB@�"��R$$X ,�R@�!B �HY �@8��H�$(�$ XP@�� � =�����aC�[�xnO��>���?3�w��S�s��ן��3y�xF]��M7y(F�R��I�7j�Vb:�]�:�(���HV�m���h�^�4Uś�.l�x�C��f]�\�Ys�n�!��z�U��݋.��Q2�B�ǎ4t��c	R��i�i�U��	���x���'�^�U"sXb�Af�*�ԫ��.e��y.�&� �iR5t�� ZQ�e�kSj�;�L[��y����8L� ��v(�r�ӏ��6�\M�om3umToRZ��)�"\�@\,<[bk�wF��C���m���e�c�H�hE%�b8v�l�������+1B�eX�c2�vp�h�Q*ܐC/m�`ce��6�xUj�4�Q�m$5�sZ�`[Q�1�i=�w2��J(�B�:c��	�C2�6�kD�%LNf*/E-قm�Z�����J�S[Y�PC�c\Ҏ��)d���\8�5���p �H1$�\vf�tF��W�2�fᬡ��R��D���W���Y�
�w�Q�h`��*�e�������'i����M��c/6�Mn�;�j������;�ĥ@=,nj�`��mEtH�PJ�f�Bi�xآ���w&�/i;?��^U���W��M� p̋�'N�bN�]Z"�]Z
(�E�=YDXm��J�PPU�C�AV(��	�r�-��(�̔չy.�\N���8D
O�NR����V�h )jr��K1-�{zmQ���N�����UyM��s��@�9��F��+*iNu�i�W�v'DE��7
̆]�{q�ֶ)lóVV����ݗl���L.�h�bαHSCm��^2���; ��N�:%�Y�νCo�_-�m��ʐ�(��.Q)�%IZ�K���ȓ��L��L�3E�aA�F��1�Ѯ9���wk#��އ@�n�v���K͈:�/f�&���X�F��3l��	����kE��rƫ��v�K�2�.��{��D�o_�Efҡ)Y��~�mnQ0-��7�(݆�Q�@a�&���h/Sѡ��wZ�����4րrݝ�fTb���X2!�)� b�h3�$�Dy w�Է�J�&�d��N;�v��9����:�!�u�Gz��6�f�
]mfV��ODuF�,��kq�Q~p�"0D}cﲾ6NQ�f�͢,Ŭ�
��0P׌�E���7B$�~y�Ե�JK-~�xH�h
�c4��6�k��l3�)��`��
 �9Z�o��EAb�n� %�HʺP�)K{M�7�e%r��o�=��T���$�ݝ(wB�6�[gX��g�X8Vۥ�9Uc�B'�Y����*�
²��l3Q�Y�Y�5K� l�h�d���t�	 j鰠p��a��i��d�(������F���db�Ā�Vw)�C5(�Z�ª�s- m�VM��w2��h$����j���R�]���u�`��n�w�UoVlۉ�i&su�V�pT'4��,Ê��e�{���Mz�T�7��]��4��a0�3`��J���BYD]�I�FQ�Л(ؠ,0bD��<�F��Dbx�Vi����M��~�V� �V�l��.:��f�+�Э�ZkX�7/.�/�z�c6�y��yE6���Ht�3�ڽ�k")��bG�[�be��Y��:j!a�OhkLK͓�K'�,:o��d�+�>B�?aT�A��?�4�|�p�	��}q�XS�?/�]OP�����S0�aʙ�Uٚ���c[B�����ձ� v��L,s��یut�6�c����{l\Í��R���>۷M��ۭ���y�s��G��㦴q3�o(�����u��(Kk�;W�t��ܛ�OO<�$�l�'����N�wa�@Kt�rY}v���x,�����1�ֈ��z���Wt�k�.���*+���m�M���v�q��W.٭�Cn��{;�8��Ϋ�r9qݮ�#�n�m���-�8���|�Λ@�v��6o���Lvu���wKۤN(��t[��=q�8�h�{�ޭ#��eൡv�z�^��T9�oRl5<����dvx���A��p󧱎Ļɤ�B:��N���V�5OT"�/m��s��;f��`4x��!�����O��TZ7n:ۡ��G3�������6H�$�˽��5[l����cj�Vw�$��utl�nN7zM���|�ѣn�݉�\S���N���&���c[�i��+�����汮��.���ѳ���j����#�\I/n'p㓴��,��J��n6�:ݦ�U��v��cP�o�]��C�5�;v`�S�o#L���ݻL� Y�'.:�m����u���M�Մ46ݞ����ŠkW�� �K��̻9�dZ�����W=�7��+&�NGx�v�z��a{n۰��|8�X�v{���!�r��f�Ul�m<&'��&�ݍTz7I��v.zX9��ö�}��.��*F�瀽F��*j�9:N�۝����CGcm����c�vw����L;<�]��k:ɶ��Ǌzݮnz[%c��N@a"v��¤N�x��|����P�u�No\m�q���½Q�N�˵���Db��b����׷i3]���o[nT�Q6%���{d����ۇ�ηV1bfzT�%Wf�v�օ�ȋ������&Ս�<�v81�����v�;O_>k�O��k���l��m��ϭ�����E�����X�*��ۘ��SS����9]����q^vT��@��5Atל��^���-��u<fmFU:�)(�ͦ�g�r�[Zv�oa;4���g�nKF�O\���z�k<��\u��θ�^� _5�Y�;z;Uv�q�հ�^��8����la�i�7���ux��v����s*�:��h�,�m\�7<�������kK�\����{:�G�=���ɀE�\&:��<X@�N��ij7��YTtkY��k�~���@�O�1��RI;�;�D	;'�8}�ׁ ������$!$;d!>�!���O�	 ��
�۶�́	��$�V�d4�!�I���@��@��n$���<B�<N$4�;C�I1$i��d	�Lx���oXN�̂ɴ��a��M��t��C<��'Ф����$�?U⋳p>:b!a�/-V8TŀM��j�&������ն�0��5�R�%{��`}�F�.����^��si+,X��:���]5�N���Y�*9�[4U�@�Z��ǆ��S4VF�yvEձv�ذ�q�v�X7���Af�� ���5��j׸�Q�X�`4cbT�0Эd	�B+"W�J�5�uS�n�F���R���2��9��l�v3���u֖Ӿ��3���O�}�`!�1�g�7qK�e�xG<n�[�b�D�F�zशP�F��'s9d=~R�m
�O&b&R���nwm�\v��rm5�O5�㪺3�;�����b8�;�G1�v�n����v�=�R�2�c:��z9Z�zS�ďb��7��8{f�v���۵ǝ�MÄ�x��R�Yx��1���3��p�\���WFC�[[�w=��z�����[qY.VŒkÙ�_C;dN���׶Ξ:�m:����Zv�cO �s���#&��`ݞR{�GQ3�:�i��PVOu֋��qÂR����H�HH�~�����V����feu��PE^N1u؜��P��v(m��+��%�n�*����ޘ-ۇ>���3�����@�E�(BE��+@	�0!+ P���6�βI!�P�y�UGIU���
����4UF,V�`�,� �����*��]Z
�T�MP`��VE`�QdȪ�DU��X����DTQF���n��*�""��EEb �V��b"�PF$b�*� ���QEQ�J¨*�o[��"��ET*�V(*�� �wlQT.��V,V*,QQQ�EADE`��Vn�"�(��PEU�Q+��#ڊ�W�*�҈�0(���"�W�(���Uw�p��Tc�+�MX�X*1��{��S�2�UTW����"�b���Y�(�zaE�R�:�Ҫ��V"�Y��K�j��Z���08ʃ�
uh*,E����*��a�(���DL��
��1�Q|J�!F(**1�]Z�ַoYy�b*�D���W����QM4DDS��Ȣ��/�b�eb�Ub%jEV�TF+Pa��
����ݨ�UX��w�� m�����ܲ�QX���E5�~n��Db��Q����S�UU�U�(��}�[�f��UN�r(��f��F �*��b""�E��w�`�r�UX�T���wUsimӪ��T�a�f�d�vg����՘ ��/�V)ݕS-_mE#G��%h���H�UV)���u�Ȯs�|�(���"�/�D\��[&"�s�5v`UTc�� �?�s��t�u���xk���<{L/��"1��	�)��'[���Y|J��V��b�F1-�X�ե~\2�ʱ*Qy�5�:e"���{�࢏���TQB�_ud���Uweb����w���=��l�X���+��R�y][����w��A�MF"*�tֶ'��Q��r�Q|J��R�6��̠�R��
)�{��O1]ݡ����Bx�㉋�>������+o��r�:o�%r�z�ƥ��_;��geoW9�X҆� �V��>�����Lw�;��-F<��ۉ�y�`��co�,�2���gt��:={�.��1E:��^��y�QY�T.�'���
 �s.�X�h(�5s��{���{q�u߹�f(֋�T���*8�V��:�γ^�2���%bL�0!�A�y��a�'w3��U1
+��\�vt�uu�;�3�_i^%���v�n�V�M�뻉Y�9�b���[�5zx�V���{�}��V ���h�Ն��Q7�%��f��E6�B���ݻt���,QbȈc&7K�`Id�6%6�E�P��Ї��Tc�j,��tYӴa��*�=�F�[Z'T�4EM���V�b���c�U�G���zёM�{��J��fXQe-Ք��&�{O}���m�rэz�,i˝f��V
�0<o)�Wm��yq�UgV�N{�i���F9㘉~B�����WJ��H����<A���;��qSC����xi�]�
{J��3�����E�-�a낑y��zi�#_L�k�T�G]]L�X�=���������:ssd*-Ѯ�u�5u���b�<I#��Z���F������]]l:�*��5�������'C�0֦+��_0��J���v}bMC�upj�,}�ه :�k�u�
*��f;�9�d�z�>���F ����p�77��M�Ӓc��X9t׷3����K�^j� �C��ck3��b0 ��_r0/�Q��Z�y�t銼˃�����#�;|e��RF+_Qj�~X«�F6>�����]��L��a��::�r��������j�Q��V����o'=�a^��k��¿ՖC�b�?����nN�f�(���r��	���<���ˎZ[��Z���7���\�J�5Ux�`�T��~�q�4� ]�����ޭ��^�+8�ݚaĮ5y��/H`��U�>�}p��V�ѭ���k�@P��C(�j��EWs�@�����1 H�?b��C����E}�(��r�'��Z@L���r]e��e:V.#�]�j�j1�����K��g��B��a�0)�	њ����O��	�[��3�9`�Hpw�Y�X�I�B�d��� 4��*M�dh��Я����I�������6F"�b0��XP D"zo&�[�1�qLCP�t����tm��Q_El�c��M��1����n��So:�~\6"�g=j�"�BQ
��M��I^�3Z��b��-C<g����>{x��B�|#k[#U��o��� ]ۖ�JyI*���0�K̭&�tك@����!G.�3"���t�	�����B����1�B�����Y<~�^i��������dŘc�L�&�+�����fR�4L(WR6���c�F�ؐ�o�!�Ń�&\K9*���!��F>�-��c\�$�i �"@�YMg�i�b`ܓ�u���(�?iܼ�wl�D��`��0��rbE��E�`��W�@��i�^�E�"���u�Y�a��g�T@��+m��*�2?Y�(`�D�MCgv��,a19tEJ�1쀸�hS�S��X��vE �R��>Դؾ���e&Bfa'�I����&b�Pb!T�ЄA���"�a�ۆ�EKMR)�ct��,U�g�
g�QT��/� vZ�$�=Q?_��v�E`��=�3M�}�$C � �z�.��QL����X�4E���n$J�����?�י��cɳ1�)�^M��:�+*���?"3W<�:��.��wΝ�ە yPD��nz��x�v�᳑{t�/8[
Ț���(�M�D�ӻV��o}q��~:$�#�#��8�~�G`(�5�ў�Q��ݾ��4������ �aD�m|��D+\��{�WO�}b7�p���'�Z��$�r��Y��|q�B[��s�>$L(��Lu5 �Œ��(Gl(�vdЍaw�݅d��5�A��kL �2���0h�X��D,��n���P��GC���n,�y@:�.����#I�2���h��>f���G0s��u����7<n��\(\�m^HB��Q�{�p���AZ+ڀ��*���,�2��,:�������<�; �裾d띯Aq�H��O���ߟ�\~�Kc�w��p~,֘;��`���`�4"���4��[�U�අAT4��ml��.�������:�8�ȁE�Z{�+[�ʵ���Ԓ�9�	k�7���C7���&�wY��`�� �7D�3�[V/���8w��|�)w���d ��
�w6�*(dTH6�ܷ�.F�
��aؓ����&�I�c�A�=��Fm$��p��7+9e*lv6���p�\���uJmέ�+�Y�`�{-s���ldEA�R� �q/���	&�'շ��1`*�u��n���X�z�����ceN!�$P��7k���@p5Lfh�t��d�R��\I@<=�(�c�T��gM6,����>q���P��� ��� Ql2�Y�z�H   �@��.NL��1`�"B����'C�m+�TNR�޽���ƾ%}��kΜ_o���@�݃9`h�$AA���d��BDV׼\��A
-}pG۵Ly�j?����
��Z�}�m�E�Q���\�wUY��l�y�z�=UZ�T���|���@��K�4e�3��0��:ӕ,��f�+T�7��?{��ُj��h��2"_C��`|�����%"�1DWv���������kW4�s*u_�N߽����~����@�%1��r��U���5T�0����ў^S�,�� D��lH��SF#�C���EF.3̯��႔�ߍu��މ�-?X��	p����.�ޘ�v"w�A�Bw�Q�b kճ�\h�FDt��2l�ge����-E$?Y�|#��`� ��8I���m����gmQ��˟��|s�x�=�::O�f<�PX1L  	�aA��&�D�<�bu�C�w%��ø����� ZlA�M��<���{맓t.�͂zV�6ڬ�мm7.p�\�n�=m�m�iӓi��SS�ߠ�8�D��DTQ��A{����$Ṅ8���O�5�U[Mu�����[�e>\H&�
���^D��SP r?��ܒ*LG����P,zW8B$p��"�u/�-�W��=��#����d��PV�:9w��$�6�g��"G�I#O�2��L�1b4! ��G�~�rb��$p����,�F�D�&0	2
0���� ���ݻ�9��cQY.��t��|<��aS/0��4�㺻��}s2/]zIi���{їb,A W���'kӽ;ٳ�ܺ���S�^���f��V�A "(6����(Y��AE��k�h�M&���̦+��:ab����2O�ӼpD��u�S�#�8 �i*�5�0��>fL��wt����sa�ĽZ�s�k�b����F6����>e�.��E���\٦�Ymv��3��8?;t{~�}��zȩ�wA�؂DEʗ�d>".L ��LW�[M>f���^4�4�͢�+o��Ԙ��8�:XlG�n��#|X�1� F�YQ�`zV	�`�mG���MEGG܁�(B_ ɀ:���Y2������
� ���"4B��7�'�$�1ǂ}U��uP����q� �C��i���@'�eQ� �5'ýJ8�"�q���0�$Ȅֵ��؉m��4��e�q��7��]|6�H�� �(,x}�KF~�1��3�����zs��z�W����ͨ�׏�E��=���0�~$R��
q�[)pʚ�&	uN�t�ф�b9�V�5�b�m�4H�  B> ��A�͏[��9w��'�;�)NA��`V�R�xv��|���0$�
���"�
Jm�]���I�Pc�aဌ$
�#]�����Λ�[?��ܝ��O��!�\�\4Cf�۹��[��X�C1y�=�H� ���Ę ��yK�6�J��c��>�ˉ�c��{Y��#���}b)+& ����Ɂk{��t�>3v��ώx�v*M��r��j<�,1xn��d��,��q%�I����A<���巋8ߦ9��
٬6����I��C/��Թ��k�ލݡ�g��H�O"0����[����\�Pc�����έL�v[�̦�+��)~��]�m�����EC�k���Vۭ��� �(c�s�J�n�+�o��� �B|d�#��U�v4�9�L���*�C�u�'�]#��.����w\�y"�XӃ�r+ż[^
�|�`��0���4����m>�YfGŚTo5�L�	�!x�¦��(�OԽ}s�jj�r�g�?c�iY
G��D(
2�L%Wq[��̛�q�0q���㜆�����-E"w ]6P��ĳ���O2���R�O���?hq�-�ve�!m�����7���d0���Y��7ُu�]Qw���EC��q����c;�s�V��Bo����B*b�H��_m]��D�&9Á0B�i#8�(^}�]5�I:T_��yT	N�Nf�7�z%ѱ~�f��R< /^e�^��l�{��T|�a�@)80�K-�Dē�3�9��/���̈��ya�;�i�V�� >�;����PCrT�x����[0�gDLqܵ�=��64��[�Yu)qU^ջvz������U���:"e��{� �x����WM9�ywp�i^c��C!�4�)�َ��p�,���^{+lˏ5��(��`KR"����Nf�&Х��LS3!q�"&��XS�ԕ�kK�@0�ɖ��O��F�<E!���3|�I�|�Y6�VZQ��{��n���>
�_��r�H�*]�bc�#T�̡ٓ^�Ɲ0{��C�!��ۛ�����7E�VA�q'4>�9�'\������!����ʋJ�q^er��:,��'J���(7�9�DG�H��gZ �UoF9���m���Art�Z��;�D��l�X�3n�ӳ�b��8�C���/pU�Ս���kl���{2t����f�lT:�NV�5�5�_���z�n��`�4����;m2�;��zx1�l�3�vݼ�u���g��8�p���v��em�6��O/;nWtm]vB9��ؓm�ܖ��q�]O<������5��[���0vW'jY1��F�-��"n]nR���ۖ����<7���3��]J0���v�8Ioc���卵�.����#l����͍(����ד:;ut�Xn:�p�n�����1vGl�zϺѦ0	F��V�f�7uݵ����������}~O��ߏ��vP0W��m�c����ǈ��ϋn���H�r��Y�s����3��j̚z�f���)P{���~�͞
[��5b�O���>�Q�-z������}�<.u��aW���/��+�=����K�Ǝ+�1���^P����bz�63��Q<����P*�Ș ��^����	�!�	1ޟ(���C��g|jlzfK��Ɏ�%x��q��]�|2�+���0�Y����.‎�짬��"O�ƚvS{�d�Rg��m9_Ӓ�
ҵ�yv�s�*Tp�jMk�#�,_r����Y�t�q>�N�j��m6�	�F�AS��n�>v����["��>�Z�m��$�B��7e�G�'+��9U�xW�͹������5��6&s���l�I�_�YV����<B�`�K�S;��6L%y�A��~ayM�����V��H�o.�7ﯗ|�ݪ��ZJ��ߔ�~sߏ�:���͗~�����0yB�O��|ہ����� �j�6>�>����ى���S=3����G����_RutЉ��>3�䔶M�yM�2vy���2��z{��2��7�����A���ɀ���i��l6 ��oTB�rf҆�E/���rk�m_52����n]9���]D(�|����,*`���,(��o�
�9��(���If	j59+ڔ���2cl�1�u<�As���kBW�Z�0�M	���Q���=	�N~_��^m� ���%e����'f���-;<ݪ�:;n�ŏ`Mt�mh��c��Ok��mn[*��?]��L�v�l4�"����;e�nc�[��H���P��C=N�x����T!���ډ�^�K��딕�+�=M@�+��h?N�f �!.�ty�n����*�3��_dU�o��^���B����$�
mCd\�dq��S�ə���_X��}��P>��Pm���qս��Z77TfUV�
W��p�0kKqC�(��q�^���q���K.MҗDr��^?����pI���+;TûZ6GqW'1�H���U��M�>e����C�Mp�E�0�bQ.%�6��	�m�7R�yrɩ�ё؉�����FU��x7o*�a����2l[b�Ӷ��;�c8�����)}���	�i9Z�5�z~44��_v�~�Tܿfܙ�.�@�;&`;y)]>K�%u}��>}kߟ��q����ݦ�����U�j��<����^u/��!(zwZe�"|�sN;�'*�C�F*��qWZMU�{Z\r�R�R_z�UƄ㜈"�)��4÷,X�'���s��c���^b��<�\d�����lBl���2�S�72���5�/�`�+���
��>-l�EQ�؆~�HŃ��X���s2�\��ɵ�G�z3=1�g#�n���ΏMlNB�D�wsr{7˞T_�p�*/^mH��^U��nن�E�ʅ:���OG����.cF���5�W�"%�A/�0J(�R�kv��K�'ot#�t���w=��d㦙3�k8�	׵�kq�VCy��gRs��ݙ#
�{�/-?~���>���Ɋ�M��u�����?,��C)l��t��xH��KWg��J$��0�LÒ;�tpTLv�[=���g���r�bHVe�{K�*.��aĕ�9�Uy�y����f�n�QK2��v�ڡ���K��29R�i(�mߣ�����y������v,�Y�q�M�D��#I��zp�~��E/Q�����x��Y�N;�o�Vr�0n�w�j0P�I�>��H��-�J���(-(����Ɲ[�K0z+���u���^�1���qˊ��U�E�z��Ɨ�÷��������j��0�ش4^C1�tr�l����WoW��T��T����ܚ?^V�]f��NL%�;sh�p�{�w�S[]��5tԫ9oo��� 5�}��;nF�]����v�;e��7�-�͹QB�啍(]]�z��<��eko.�w&�7k;oU� 
7htur:��3�-�{y�V�&��i�sU�&��v?C��>���3��2�mD����V1��dИ�c��!�Pfo�P��{��s��؍��������~�<O��s���Nh���Ї�a�)�R-��׼r�X�E�3�g��wFi%�U�`�/��-F��i�(�Ϯ������q�W�:>y�#�o�g��\�[��I]J����[��`��X>ذyS��# zI��m���e�\c��s�V;�]WvlC��m��c�ʌ�RD&�ʢI$Ų�a�L*j�/��)�"�ʉȳ�J�g��&�ʌl��(@�fb��m3C�dɚݘ�k#�ɼF�/hJ�^�f5F`�����0Ng8���<r�Z��tv��]p��Z;��;��u������U��6��&�;4Ka�@e�����J����:��vڍ�Όp��jy�s�Sd[{�^'w�!ٵ��Z���3
h܄�9�Wca.$|�����b3-��{*dp�&:_�:��Us�`�P�%4A' 6�6��}��� %\�*2��¶������e(�03�q@Pimtt�a����j�:}�3���GU�]��V1�+3F)�w����w{F�T���
�Kb�:�`�c�'wj3*
�q�X��ɺ�2X����/|8�"�H�t�@�i��d_x�"�TG	;��*�qhB�����c��u�����W���i8�tn�y2'Ԡ�
�Ǳw���� �p����:��D����E�2�?���}��ϻ�#w��]�nB�ۺ^~�*���,t�+� [m~t�4CM5��˽��*v�s��k0��YNmV}p/����o��_X�g՝5(�|介3F[��}��q8u�YJ�?y$�vwN�Pcl�Vկ)����*����=d|�)��|Ȑ�S��i����K��0�l6�A���Z�3��TF�j�jp��8*�%�s�/�������m�Z��{q]W\ñ{M�(�j���8�`6�q���e�=1B�ƞ�����[hǙ�^1�&>�Θ{<��t���zN�Q��. hΨ�a
�Ր�d�hI����݇,.N���1t��ڊ|��=hۦ�{[�wX���r�gm�M���.�I"g<)LR���/N�>̿"X_��
-HhҼK��N�Ӓ$}e+�	14�L��׼e\�K=�|iMy��%�#����z��6��3���e �`��%�����b��]��A2<J�ޔ�Է��Q72l�Q�ʗ�[6�p��_wf���z��%����}n��"�zU�p�=k-�~>/�e�7o���U}��H��ݻ���_/=o�싒�P�pۀ�i�BYup�L�K�[�W>*7���Ç�c^�E�/�j��I�<y�0��X�Y�z�:�Y�ICfL��Ŝ5�<j���B�z��֥'�#"��7���p�u�̭��@DO_+d�ٗ���gf����50DLC@�!�h{��\�8���;s�2�ey��'$�ѽ.D�&���5mwѨ��ݏz��n�5Mb��fV0r�H�5TqG�jr{ηʜ{���,���9���s
~X0���-'����r��_2$��,[`�G]@�@Pl6�l6�u�㓍K�����M����G}�;Ⱦ�xyMp)U�d���g�s��Xj�\�P�!&A�o.x����^�X7g�z ���֩�xP����]߄�f�}u!uį3$���"�M�ӷ4�����R��E�R�l��,X=���;���n�p���cO�f_D�p�ٕ�̳&�\��n�Wm���I�,�}�7e���AP��f�3�ub,ٺU�.u�2�ۂ��2^���z�Y�zu�c�㻶u��'��״�esc����U��#�Q��4�5�@#9�FAH�����tX��󑻁1���ɹ�sŴ)me�9��;���u�C9�7�1�-1�xˊ�5�]k�cJ�c!�[�v�[v]؂H���c�%Ǉ�ny�.1�X=�0sw]�9�u�zyϋ��xc�q�eCYp�zx8��h�=v�l�];�8�i���iǷ%�s��pm�� ������
�������]��jw^�@9�b�N�s��n{t1N<�M����]�;Z�e���l�k1�9�8݋�9�.A�n���_Ƿ{��Ͼw�����������kQ��%Á$�u��kyѮ㝱���֝�W�=i݃�������<В;�`��[������iό�t�����V$�,A/6MR����*j-F!eZ�q�}��$�ǄOf��;�c8��ﺀŀ=��.�\�v��˼y{�'���qvX�C"�0T����Ț���P�()�7L���Z4[J�`��l���^�*���"�.���q�#��.h�lE���B[I�]`����9wv�K5���Y�E�e_3�l63�
n	]e��j\iZ��;����r*)Q�����?���_}�9�Fy3�y�g�?}�?JP~��Z���j�n�KJ�&B�q��.���I��so�}}��ױ��Rd�K��w��Hjx���c���NZ�.\knC��}�;�g�p�{���������K�����!�t������Df�9(ŚW�̬��q2�Z��x!̫S�ū%En9뚛9��3���@p�����墩AY2Im���%�#On����q,���H�w.�LT�o��� ��9�R�|��_[�ߴ�{]���c+w5h�w��-Dia��.���tI��v���%*���ͭ�o�T¦_��!�F�����=�7��
��	�(�Ϳ=ɮ���[:�j
ŷ̚���M3�S&V�E_v�V��H�V�@ie��t27���nٷ[d᱒�N�=ձ�J�ۜq�⧲W/��gtr���=Xݝ�܁��-��8���n�����z�~ڙU8�MS���{����2�'}鞊^¶��"���wt�U�b���o�=���4��و����Q�3'��˷��U���1;� �� ���Ie	��Ы��̺��uW�bv��ҭ䇗{�q��|��Q��m�Ǒe�U��4�w�P�����n;}�����KɅ�ݯ[9?BwjI6.Ru)W$��{�LA�z����&֎�vJ�Oo�S�M@��"=��$S��ŧ�+�R��3�4�Ѳ���x�n�c��lco�T�=e�;f1���qpH5�{�sU��V´�ng>��E�nH����{ʍ�����X?��]]�=�Moӻ,:D$��J�V�j&$�8�Pkn~�{�N]�����PCۀUti�WNL>�&�V�9/q���hb�I\�.���;��Q݃�)_}L��%�c/�ٌ��ϗX�e��Y�NȰ=��ѪS~z�{çFK*���ȳ���"�D������H�	Bim�-^P�TLȺZ,ڙ�JW'&�FH���Hם��5��#d$a�V,�Ԁ���}��f�S����S�o����^Ա�\�!:�ȫ��U啞.p����F�k��k¤�|vR�Ճ"]�<c�)7I��,����&g��k�VwjG����ͲQ]u�uZq�]mv��ڂ{�z�]N6$d�c�,�֙���ٜ,fE\���}�wQ�F�ʖv�_F^l��*��<��X�/kι3G�H��"�w�#U�+����ײ���1���f��9=�r��YgԚe�_�� R%�Za�FA
,"O=�!&���ɀoa=�Ce�/kG!B���e��4g�6$b��(�F߷�2z�{���q=���N�Q6�0�f�������V��K��J�Q[�����p�2}�FL���)�i$�m�(���6�ٵ��bq���Y����cq~&�Ǧ8p���.S�h�G|�Y������0`f�/6A�aܙY�·u3��j�v��2,����'�ԣaڐ�r$
��u�ʷs7�����F��0C�Z&��b�"q�����Q��J� �{k�}�3X&Q�X*��X0Qd��,���n�aSc�rw{�؄��j.��%�*�#.�������Ǐ�`4���g��#͌���}�tq4�����O\C��fޕ��e��l��7aY��w��l6�4��c۴��h2y݇��,FcQė�U�#r���]("4}#����M��q���w��3�ʝ&�}^Q��s����ul�����`F�e9���Wwr&aM���m]�ջN���z���W��n�0�� �g��'�`��M̴����.�������M�ٸ��qכ$�r������+1w.�v�8�JYB��������;3���&��\=�e1��U5y�PHc�[�[��=;�{�W	��f��%ʨn�j7
b *B�����0���wIY�Y>w:Gg:ͥ�Y��'�-��q�5c�)j�;����۹���(S��X��8<�w��7a�Qwq.̈́g���R�!�$�Υ���Hl���o��	�َ���0�����# ؆�0�H�O��;�un����=�v���YE�r��bɋ\7n�v��:n�Z�t�R����Џ>��0�_=�ٌ%�o�lT��O�͋rs�^�UY�Z�ۉ��y�N�U�Rs�tӉ�	��O���J�͸Ή�^QB,N�U�?a����d\�B�� (��ED2�$�0�k>ك��.n̯R�9nl#Y�<ҦyH������ �Yh�U\�4�q�7�K�歡 �pTsc��R`vLP�ő������
H�I��`�Fķ�[ʫwv��s��.J}fš�`cM#:h2Z�A"�c��Jݫ�J�^��l�?n
B��#��蛘����-6�t3�AQvWTS��}l��bQ3sp��0!'�W�u�9���l4oIv����T.�l�����[�ݓ��w�ߕw1�߇���rM��Y�幕wQ'0����Q7F�&�V��^{�#�~���3*c�ﵽ���9�S��Yӷ^#�t=���÷�<�x'c�;��>�$�O��c��,zzM�)�����v�7�Mx��y�7�`��~������<`��%BM�m�y���T������Ng�I�+&��8�71ӄV�A6�9���`;�OR�P�!=����g�X��{&�c�p����a���E�E�8V��}�'K&����Kɿ 5��ͬ�V�,E�i:s<fǆ��l�DlƳ�/b�cnJf�pu]��nkb�S�vBrs6����u��_4ᢚc��U��Z,=E=��K��3&Ȉ���^��X՗R������xV��R�Y�7WQ��R��M��"��"W��+e�1]!��1�Z;}o����p��=����P�����ޠ}Q��ݎ�N�|����ܭ,4�PB3g_�y�;����;�ӹ�-ܡoPkk��L4���H�{���3H��tI|����t�q��~O+��(X��U�c�+;�6}Y�"�gcA�ʃ}�",�A�&�")S,�����2���[{�a��g���NoĀ�0�fe�YP�'ck�E����&e � 
��{`�S��+���&�U�:Tt}�˙ū��`�\����8Z�c����$�e���7}�+')X�f
Ϟm�M�1��~����|�����S���z��:�b�y<��A�*���N�+i��`�c�H`X�S��z&��|#�2�����-�WS)b91�~���@VH,��M�a�N=>��l'��{�Xs
�Qx2�m��F�9���)��b	�*�x�]�HEZ��ۂ7�kn�Tf���p�6��O:��z1�bB���3�?����r�cc7�u�vՠ�\�w�G���<86���l�3����0������9�#7ɛ.үcIõK����$��Q2�1U7"��R~*���}�~�5���9vA�F��&Y��5	e��v�+�Oj�f*�:om�C����Ρ{�̻ˍ�pjzٔ�,wI��ie>��I_>f�'�{��d͌�h�F��0��+B���/��r�݇���.+��6W-�����nu�0;�A��҃v��㗭���K���Ϙq\Eq�e�a׌G�6㭃I�N���J�MOgn�yb���`�f�(�s�E�7a��;p����s2h�f��<gs��h8�]��y�9��]�>�ne�ru�Mq����c��|������[i����s��^$ç,s ��lv� �7'<Ic%�Xb�ls�#m�f�y���&�8������|^�='�s�ױn:�;V����ݵ��׶����϶�Uu�v�yq$KB��m졕�[���,g]gw������o�glj�#sq��������8�}~�3J���|7�������b��<�R�C���<���p*�9�B�y��C�,�@P�H������9[y���:�۞��	�s��s���5��q�έY�zV�uz�ﶫ=p��I'r�b��鵭{�z��X�j��%x�;w76we��Y��pus���$�c��jh�и|Ɇ�B�ၵ>0�&(�=$o+����v���f,.�{c�h!9[��3Wu��x=%�7%���=g��p�������`��������5?b�1��;3�P".�m��� �e�h��Aw�yM�.���O�N�����k�'O�d�%ІБbۘ{W8o���3h`��2��i�1���w�-���]�0�4+`��s���$��]+=��7���qn�R��k�����M�,�p�I'*�Ul�':�w{�o�m�Cu�Z!ޅ�p���`�(w�4_�D�L�,��<�z7��*@ټ�
'���/�׍����3��o(l��cR����|��^��2�t�˖���)��*���u��7n��ݫ�znq�-ۛӎ�[�Df�3�v�nS&d��������7��O��ǳ#@Js3�f��bB�(\i�J��bn+'T��!w5p�ӽ�ԩ$Ul���g�,��ѫg���&��D��6@P
�(6�M2��&��[{��f}��!��BV]���l佖���9���
����+w磅^���oV����ݪ;vwt�Ց���;ov�b���V��}���T�@�u^��9=WQh�\E�������	6v�B2�\x�z:ǳ@eܬW°�N��	���$m��Kt��z�|
��.�K�o"B�0�h���/'+m�=u\�^��=錪<#�쎬8 �h�C�(8l����kd�+��y�~�1X=q}y.�m����Ƶ ���[���>fngx\Ӈ^�s�;&W4�@%�K.�G7j]����8��w[JS��
xH�w��_�B=D��N��٠[o��K�9��6�w�<�{ۂ3�J���恬T��ݼ���A�*ʛ}�1��U��*	HM�z^�TF�S��}8��V.�@_'֔^^��Z"�8nƢ�2!6t{]u�Amm�x}'\N㫬�}b�;S�\������ex�؞���S�%�����Q)�x��2�p^`�,Z�-dF�^nf����ڞ�YmE\�A����1z���� }b�4����9�E�������1��Y�+;!ռ!R������6Iặ~����o�>o���׼7hZ�W���g��'�v̩�:�7'g�k���>eMˀ�<����;Se	�vw����yN}3	?)��7�����*�@�S����>)[9Q�� ��!��I���m_������;���7c۬��8�`�>��9 ��l�}�4�uK���c��R&*v0J�J��KEv·���2눨��m�5�%`~�nȾ�XC[�/���N]l�¶���
���.gon)Mnej�v�6��+i�C37.<FliM�U�;z�)^[6�N���;����ӌs/�%>T:��k���棪�Ve�����9Sf��G/p�]��/^VN�j�dXwu���N�c	�"oe���#��&�x���j�.�������
�f�z����P�f,p��[���2�r��J�f�
�T�n̦6bk��٪O����f,hZ�=�=�[�����ӕ��QW%�٫M�5������J3������˨�Q���.�n�}��S%����r潗�~��<@�U�%�j��ǵeA��ZH*@�>���wAS�.�R����mPW�g6Ի��7t�v�Y�}�n���Y�J���nؾ�/Edi��Q�t�޾��W��s�������:إ<��Y�5`k 4C� $�I޺s��b�8b��^tq`�\���Ǣ�F�ڒ)��=��a��E]L�1��7�/ޛ��1*���-ߢ��#I���I�]����3���}N���I�="�;��y�8=��x�7�6w$s��ҩ���Ғ�P#;̨L0�2RA�)�M���a:����,�q��ܳda�邳���J+��X���_�����;/�ҳ�]�jn?��>֌{C��̝¶;��`'d�
��t�*�>�Y7c���ݯ0<7a`)D6�6j	M"���8�/�M�uy�}�ѓ���dگ#�l�F�{}���B3�+��!l�v
�bN%��ȩ�����7�=Ʌ�=���C"I6�QfȘ�!�F\�w��kxid$��e�k�r.��\�n�%�����ԡ[�$����W���;I���k-��q���jY�ݒ��Z��iS�3�'DŖ2�xj��z������Vm����|��m��ն���f\߶l��\a��l�� "��J��d����+.f����݌\9 r�*>�/tU��SYWtsp�u�F�q��T\N��7�����w���C����E<�˻�;�}�|U�2_\��^�&V��٘.A�	C-]�]�b�U]\p�cp��Wk����n-<�7�N�u]=��\՚�~K���;����4�l��=L��v֝8{���C_�xmڪ�ܴj��vL��gukQ�*'yB�#�K���$��f��cK�W�3��]�x;��RF�֞�v�,d��
d�r�fdO���^9�E[�ͳ����X�N>tG�-�?��O��͊�Ǣ��׽g�?`�����7ё����4����}��������if}�,f�(�}-y^�y2$� ��͠�7uT��rb��2�Y��u�^٭�\v�j��m��,���~�t����C�l��G��f`Oe�v����{}�8�/W9
<�ZwR��U �ױ��pyd�sKM�}�w���G�[\7m��AS���&}>;�B�y��y�"jB����7v4�O�r=惓���p��c�r��F�צ/�q�Q���W_K#V�/a�D�"��Lc�ڵ����wv8^�wP�����y�e� �A�e@	�7��N��j��}���lY�	qVE���^�{�p]�FRe��flE��9{w:Wq��i�SL���b�o���hJ���W�B�%r���.SbX�oܢU8a,#CA���R��W*�j����D/���;�Y=[4~��ǋc��(��YS�jfY]Bu�hb�O����[�93p6sk��o���Q��,�L�n2V/�R�U�ջ��73?X�GP�M���#}q6�C8��w��� ���z���a�}x�Wb�*Wm9�ܒ�r�`ةy�	5ث6���8�=����%&
F(�4�^��-�ͩu��=n����w%�p==�>u��;a��6���l�<��(����q�9�5�xڷ��k�6u�En��֎LT���48;3�ntq��m����N��*s������0ƃ��tpi�Q�D��xZ8��Xv��6��k��2�cF��ki<�=�z����2�ksm�#�BIn^z;.�ۄ,�l�=�;lqq��_�����i�T��lV�?&1����f{`��٩;?���������}�����틔u���v@جα/�-s�%���9CŶ��#H�S��n3GU�s�/�1��D���4@�m�TL\^�����o4��secB�^oNQ����]Z_��v�O�p�7���2.�-m p����vº��V�S&Q?&	"\7�O�2e2�ٛ�ҏ�"�o{b�R���_,j�ؖ�ׅr�F0M�,��w�q�����7�e7~�CL��r�VG�6�Z����FR������T����N_�wws1�5��^�Ã3������x��^o,~r�ڹ�E�O�g��o���ypPs9Q+/ԉ����\�F4WB���3�9{���E[�Ns�hL�=�]g���R����v̂�Ɩl��S�~m��I���!�m��A��6���J��q>�+�����	�m��X�Ĩ����cQo=Z��'�EO�xR�����Ө�;/����	Ŷİ�+~�S��2���=�o�Tu�VT��9���4�	��R-|Z ���/u�Nzn�>'mM!pd��y�ޛp��B8R�&Kh�[�`3��� =J���^��s�ײ�hbuS��Gb9'�ǽ�IY��ԍ�*d���XGƧ+Ő� &�i0g��n6��C0�BAi9�yG3��nk���C�z{BY̶�W[X�n�	�#H
h(-�1�خ�#7�uD�����U���u7�O6�G\ݾ5��wj��s���隧R�d����͟Vӵ��¯$:�+�b	y�>p�^�Y�D���ɆIhC��;�^�bc���ߧb��⑷�zM�~3/�ʶd�@��k��Mg�{ӝ��߉�c̃3]�SWUb*`������_�J��~݇O���b�Y=��<=��^7�|gl��ݰ���$4�4@*%2h���u>�7}�j셕>����G��VW��������X�A��SƏ%u��'*�`�����ز]˫���w�bɘ�����c&Y�y�\fQ8W.#n�ֲ���Q�V�m����XL�@4!�$	�����88M����Ӻ^
�mu�]f
�L�~ƴ*S�H��J���il����-�rv�X�*f�bЙx�W":ۭ.��}0��}5����o#�~���⃮���?��^�r�*�~���-��ϊ~�>��ϦI�MA9��ܜ�˷)��z�6ins~�ry�;��l&���{ُ��-�s�2�҉��Dl�w�Β1^#togw爥�]��Fy��`*����ݱ�iƘ�p{����ֵ9�c�z��D��M�s�&cj�k���_��}o��}~��o�q�.U��B�l�*�KȪ5��A�F�l�^����v���^����v�e����f���M��?j�_��'��.-����~{.s�à�����IO�b	I��c�Uc����n�cf�\T�d���੃f���C|֭��o�o3�)�v�&��+�5y���kFY���zF�Գ5�f_J�g2��*�V^o19h�噪�����{���l��,�z�.*8op��/vOT������9��b2�[����򫑀^Ԓ�ν��b��5f�$4r�]�rlC������냭�ٕ����J�H���6�fS��4��O����n*Z9�M�hڛ���0L�t�3xJ{8�*QW-������?��n�>mC�K����%`��tu^��v�z@btӵ��Im��u��ʄ���Y�[c�C7�W�Dik*M�;��,Y���}�Y;?�xo=�o԰�E5���!���u����˴��7�d�>i	^���=_H���� �!0Bn
�;�����/(�kr��>R%v^t��٨���ц3�k,"6R��d�����{�����������u�^M"學o��nsG&��[ms�;6&���ʨ���͢�_�$�
��V��y���ݲ�uyX���N����W�c�`Q�iUN+�Q����NŃ�Z�}l���^�FH�7�g]L�3��X�v]���/vUޱ���'T�yF�Z�Qs]g�3K�չ&��ؗ/73�^��ĔSѵ�q�"�Uh�࣮.]�ɤ�@2Ra�6	�L�޷� �[g½KAŐ�2�,��h�깆�ܭ��<�6�U��>���(��w��in�M{�s<b��r�x��p7��	�X%F
M���{iz���2��e������9���3
�8�X���N����p�n�ܺȴ�+S��yͭ�V_<��yZ6�tm�Uk���o�k�k�m Q���)#m�����|8W��B���`�A8L&a�V�{�Oʾ��-�eg���Ώ\��ꬹ�������Y������9僜���ʹ�	.p��z�/gCj�}~s����Q��|}���ϝ�U�.��wz:.��l7C!6>I8+�8"���3��*�W�����ay*�e�:�S8�C}j�,��M��1�1�B�p�vo5�$k������D�jv�F�p�2�'��w��8��޼P�"��� �9��â(Z��M�\d���ӉP��!�_c*Y�'����lk���;Z����1��Fd��Es52w �ux�P�ػ8g�ֱ�s��UNv�T.�9��9�z�Դ�N����^Q�� QN�!�C��=��u����s�=����ϐַd����Рp���۞��^5	��ZIC�6�U㶾ث~�C�h��󨑙�m�^�s����ttt�G�Hv��Q��C�T�MG��`�8�̕�ٺ�FWWC�g�d�����E[v��sr�,��6!�SC!��<�8Ыd_�ϳ�51����9́@c�č\�'ko�K�,�u��FW�} Oz6�V�ٕ�ѳ�q�����o��Y==�lM��{E�?L���+�rc�[ 8�K� 2�a��U��t�i����˼(��w��.T�ڟ����/8l�0N�Ɲk��t�*�g-���l^VZ�].%\��B�7���yd��\�4�]�m�V���=�^�j�CII��,���ʦ\?f�cVGBO^�JEo�V8�_�m����N�n�ܚ�d�p6}��^��,�b�U�9�=	Nv�L��d��xU�5Ș�čV1��@_@�wH��,�U:��ie�<�b��ӑM���w4��P�e��G�#׻���f�:ţ�:T3����Բ
��ٍ�����S(��e�p��vg�v���~�yʒ��taB�~3��9��;�{�]��?�C���b���*��JS�$������>�~�@�_�s������A�`H�I "�I���Vx��˛�CI�H� �� �[au��BR@��"�(���5$����I4;�	� ?���$!���@�kBt��6� ��	%d ��>YvB���m{g����a�D�(v�I�3�� R�`@��ԓ���_�_��=��_^��_!�W��*k�[�}|<|�u�~����=����ß`H2@o�P�"~9x����߂�t��)�q�N?��/DwLx�����j/3���V ���$��#�1@�7� UE�DI�t��@�$��l�_����'�ӂt�kV��PY�BT�J����� �5c8Q<���
�ڿb=pz�6m�H��fw'���	�L����_�)�?��Y�}�`IW�J��^Y��۠��:9��~ ֔ı�ߺ~��������������}d��R�N�e�Y�ڽ�֬��$݋�]�{z.��F�̺@��
�ܚ	Zz5k���Cx��9�n�J	nmJ��r��T�j�BnaV?�vhZ��%���ui�N�Ê�h�fmӦ�����Y4���t�+g�ǻ�	��+m�b3�^Q���G��@�w�3&-II�~03��n^��%[O��Zo&lt�oE�n��m��kY�Ż2A4���C�~��s�>�@�Y	 2 J�@�eB� )	,�� ��D� @"@�!� � ��$�5��I-�=r����mS_��87�?a���@�HI�³m`������C�u=�?��~��`hs$���P	�߀������d_�a �f�l�� ��hv�L42gzvW�|��0�Y/�O!�&̅�O��R�ۨ��<`P���a�,��uD�]��p���T\z`"8/����������f-n�.�`�+ۗ �9*(+	� �S�<�Lz
޸��I@�<Ç�d,��4��� $��_��a��b��j3�l��HL��)7?WXa'�@�L�&��E�,,���p	�s�95��$����B�O�è�8I,6g��W��=ghWh����Cս�(gDQ�L�>j��{_���i�?i:j�%(ڙ��2 : i$��c�b$��Ace��9�	đ�t��"@�
���^�����<K��q�M���c�0@@T������آGA4����y�����d�0����nB�%e��[�� ����Q᫊��(]�4� @�u~�}!�0Gq��>��D$%X�A��͛_kx��{�	߅��d�&�1�\`*����.�e��I(j���;��T]#�
�S|J}Lq`I=��ˠ�����TA��ɫ	 p��f�O�]��BB``�|