BZh91AY&SY*hN� ߀Px����߰����P�\ۺ�+VԄ��I@	�@hSO@����C ژ����L�L1 0 ��Ji��L�SF�44 �4�& �4d40	�10� S��I��D� �� ���Q� ThD�BVB!>í~�#�*č����}��;&XA��`s �����3u���/a#K�V�(�]��n��ķr�Zs�=�1�f��h[Z�7���K��t(����vlP���h��{�f8xG"��8����I
���:7�c�^n'~���d�S��w%�HE���#-�Ce��8�r�sri�E�"bd0�B�5gke�m+x�I�V(�"F�LY�T��k��Y�� �� �K{�X������«��kZ��T	i�Xrq�.�AQ��S�I�p�
H���3�T�#*
v;M^]ؙTX,E��*�B��*�r�H�D��ޯL��uFbT8�n�^׼WÕ5��6���j3�u��y�ieo�q�N^�xب��J�0DI_���[�@l��^3ió3���8�drKL�� r�!L.G��Sڄ0l2DXBnh�H�[,l�a��s�6&L�
�)k8;�Y:�d�}����n�U,2p����|�};��RuO𚽴j�!�p�7��`HCy>G��A��@�j	���ߋq����s�q$x�|�?�6d�B�Q��Hiv�YW~�mh�'��k\�tWf_�r$��A">�G���ޚ������&$��>n�
)7'f��߀���EL���Բ�W�������!�H�;���l��`�4xj&�J5ZKqБPu�dϬHHDK^ɘ��>q�.d�֪����a:�tD�:CVt��Jo�Иr䄊P�H%¡Ok���{������4:fO:I�sݠ����9�cz"J�&K!Y�HE�̘k%g�<�M�s��"�$�c���Ƴ��	> H�]��{
������$���BYɬSS%�i�<���2x���j=�3���PX�� m�B!w���L���T�)���L�vGIP!�ׇ�a�e��2�F�Y"[�Z@�'���<���j�|�.�\=*�͇�@���A��l9�R���!��Z �8F�i�l�8�R�P�n+������̖�c2�0�/!> ��;s��i/Tf2�I:I��jqL��T�l(_�$U�C��
4L�eFV@OB�.[��}��|���L."�UPi�a�V����d��YT�#f[��1$"�du�$b^�剘��@̙����?��H�
M	ޠ