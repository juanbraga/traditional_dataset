BZh91AY&SY�֯� �_�Px���������P�8� 1�ML� I�2�44���=�=T��F�C���42S�jJ� L LF   !!"C�6����   dɓ��&	�F�!�E!#�O)����G� �bzA4åE*�I��HPlI#���O�Ƣp)�Q ���#�����k�!9�N�-���x��
��b��F~$�}_������ٚ�v��G"(�6ds�i���Y�*v���é2�eW�KJN҃���=&������qf�
�[�kmݱq��QD
��5�6���q���d̈́9&�bG�nY�>s{!�����d�.Ù��kt�4h`u;ڲƎ�3[� ᷧ���ʗ�������� \p�	#r2R4C:�g���b���">�e�S-&ն$#���lc�)���5��%���!�L�<4
ЁL��l�0v8�ru�H���q�[d�'H鴬�gRa���U�;8`�*�m�� ³D,�h"P�i�B�f�3��ڋQ:k�TQ{tҊ���w�*軴I�KD=;��'��dF���J1��-Z��,�Q�Tk�U�Q��j�M5�@f��7��K}���w/{�i�%��K�z@�@QE��k���q$~�4��W�^�]z��`��rՆY��U$,��c��*��zds�����6�nL�32N;�C;.���P�0�O��������f�����_?o��/����(~�O�w�����o���]]hB&���8��ci���4����`o*9�;�bĐ����[�V�oҬ|I�4�"�Q	'��w�qŬ�rQg�%7Y��nq�y�E��?�6���s�C7r]nRL���|!��E=-�T)�|��ؘ���+zg�Ѕ������b(��u`z#�qR,����5�	z�Iz�oϱ^aM6W�����\��n�˘ĂE�J�/&�7C&��^��j�D�-d���waSi�+oG��8Ծ[���!E�H�`����8���ya9�u�4�.�q|䪑�Q6�0ߒ�+5�h(�:� �Q��1���U�I$@֢��d.�C6Rq3�(��-�_'.b�*�bSX<�!J��6i82�W�Q4�'!Xq�6�G��{l���i�x�^��8��Y&5����l�(��?��N$j5�܁�B�:��E�畆�l9ZR�c�!���RD"��w���fM���N�Bg3QH�IM���0�X]V���X��6I��H�t^�j-W�9�o�wR$1�B�29E,Q�W���ȷj����c�~hB/f^�%+}yP��v�d�+�Ɐ�.�p�!'�_