BZh91AY&SYU �� 	߀py���������`�|�g<�]��
 	M�#MG���j=&�h�   ��	���H � h    ᦙ�&�`L#��i�����)���4�� @  DMCR�j�i�FC�h1=G�E4Ѧ��i��L��&��m ���0+Hw@s���#@	��=�4�R������`[D�� �!�+2=�P�o�X�h1��x��n�o�PiQR�iDD屦�5L*%'�8�[+��9�:װ����jt�Mw��G��`n �n�7Be�	R컹�͘�6O�xw�J��I��a?���5�M��)L��]���)�E,�
� ֿ'�<�f&(��.��n�8� �BP�P��Za�"��Lic�d$
�21^%AP�CR���+J�')),,B�������v��R��p$�L"4��R��%�&m`[T�NH),œYL�"p\�+�#��	!�»8�p�jQ�4����Ɣ��%b
颡a)z(\��L-h�=ά7^���b�\.�ޥ�e��WN��kU�ϫ}�Ax�2̬cZ�PLJ�1I)ةV�!(5�*�D؛����t`�̉���87����M�(h�h��\���8ie�n��*�B�cT�r��h2&Q��Nr��ME��)��iy��h�1QH��'��%���6�k��"j�B��:v�q���f3lET�2�J��2��=���� �I�F	H�
��δ�i+ѐ�K�k���bL5��t�@׸�$�-
�+���O��c!�IHR��u_����;KFZ�h�x�撂��C��Y�n)�u��}�0&2��J��̣��rQC�8=��bQ��àk1�$��2J󠘮��{r�A ���W|���$��A�IR
}k���[���s�H���s�+�!4��)Ӿ;{���9^�Ui����TzJ��A�@�����dk�׸t���� �o��\@L�܋Wˢ/�o<�n�+z/}���⠙5
����F]d�G-3��RR�_Sb�!U�P�4����*@�D��;w��gi5�"D������6�[qS�8�
e�L����u�b�Gi���6r��Ǉy{v(`T�^�X�۟A���{��bQ�$����^�D����$Ӝ�v�>V����� j8�*��D���R<K���^Ʒ�̀r���Z��:56d�$bT�m++�|�.S�Q	+�钌JA�|6����DM�j0R�!KMlz�R��.��ᕆ���+�'Q��Ƽ���v�=�Wb�-��9>F�`:ݐ���j�T����nu+"W�z�W`q�D�YK.)i��x��u���.- �BK2pÁ]���o1���ti�[��&�L��zl9��,k/�DK��p*����� �Z㼺��ۯѦ�Nܴ�'M��d��{Z�W� ]��d��C~�>m�D'y�Woٖ�� �� �������ܑN$@$� 