BZh91AY&SY��~ e߀py����߰����`>���i�����Ph�В�oJm�4��=OPP�L� � J�Ҟ��&� 2�@ ��=D���=@      i!D�6"2�ɑ��A��  0�HB=L�=L�  � h D�hF�'�����&OOS�OP�z�h�jhdP�0�z�օY�T$ �}��$��uI����?H8�� �"i ��*���]dQ�#�¡4�<����.}m��=���"q��$���� ��붲Sj	����Ip�􊉔�ь%5ꜨN������<!B�6Y]�\Q�x�Ԋ��#�d<��GeR�j}[^��L޵�K�S�����v\7�W�S��%�k�7��:�vv^�&6~:���� C8�&��C선�-��Z��]r�ݟW��s̈�"���>�c�^4[��t��]�d�s󣴁���;����;��U�z���V{�e|S8+4F`���\��>(B����k30B�:�a����._�=H��@�
'D��4\"X��e�>qC�Y�H�9<t@�mof]�t�r�T� dp��P�-k1�E֛Jq��UW-R�R�<)��rq��l�vZ�V���Y"�e\�c��$�sA�V�fϭ�4Y��}{�S=R3d;;�a}�Y8X�h�.^��+F>�0��<`���P���6"�R+`�H���(��JZm� 1�+@@@Z��^��v�ʲ����ۊ�"��`�m� ��z%�[H������.�鐷����)�w!m�N2����t3���X`��*�ՙm5o`��dZ��$z)�L��M�qD�v��I�����=0��#�b�1�Ң[�b�Y��Wi���Ω����eo����<$�H&q��AA�C?�K{�� /ëYv�/\-Z`T'�%���dF�pp�%�%AH � �o�$������ܗ��0T��[X_���,+-��(����Ф�!�6^�|k�|�ׯ�rݩ�¦Ԕ<��D
]��8����37���a�\Ⱦ�i�dD����	�8eؑ�������3���!^�~��4��%��u����]֒Mp7kǆ�I2�e싌�"�O��ǳ[W��$��[y)�[.�
��R��06q�~���2~���Ļ	17E+1vQ�bُ׷X���rS�o,w� &���ym�OL������il!A'��&��Id��$p*T�AA w�,���U�0̱�)�;��D|���R��Z d����{A��V� ��GD0S
�",,p��)���~�CS�C�K
�t,��y��4蘧�O����S�%V�&�Sa��C���w�E�x�K��M����lw���}�4A�넌'�G�şJ���LS�i�:��@�9Z� ����=�W}')�f���P0��%\��ԃs~a5����a1(�.�d\� �����E�:˭ꑳ(}����.�2qd����%XbՒ�#��Pi.3�8��R���y���Y�=��ƀSNM���ɚ����>u֥�nhoKT����H/!Ȥ�x���hDA����
B҅�|��u�A�ۆ6��?3.{u��;=w֧ۚ��.6KQ���_���~�㝓�j�)�t�e�`�sN�f��$��/�ߐb�դ�q8	�M���+�&�zo�(�d��oמ��˖�M�M\5�����C�y�ۼ�O��&��nAN�EKKRI6�ڤម�>���(g�����T!�0C�bx�_�rE8P���~