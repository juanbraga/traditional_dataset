BZh91AY&SY�r��(_�py����߰����`��|H�   
  P   �|�U*��"*T�QT�
��D�r  ]�i�j�P�����T�m,P>���ޜ�۬����^�:{�48��iB'��親�����(�6s�N�l�uR'8�xX�(z�@�X(�t�@<ǣ�/rp@��4A���ޠU�jpPi�t��4h:[��@��G�tP4a����t���T��� S��a��t�t�AP<�AA�˃A@���(�A��*��U*�֯  =ܸ: :C�W
 u{:t�/V����h7`����A �*@ 5O�T�CM4h4 ��2FM4j��bi(���0��0 �  OF���T&h ��  �C ��TM
�L0� &��  �I%*mOP ��OP�h��"���O!4�zM=OS1��-F�^�k�襳0��B
�|�$�ga&��	,$ �>��h�	$ }����'���g�����$��³���-VϷP$�60��C�l^�M�M$!!ZV�ۧ^�r�rx�WF �^��	6!Zā�!�(
 $*��CH�$�$� B$	*H@4����T M$�BEB)�"�I R@!	1 $� ��HP!
��E$��C��%�>�$�\�d荎��ʆa����A"q酒�1!U}�u�+���&a,��dŸYRŮy+N�u�W���3�L�����(p�X�"M� ��r�RQ��n���{12��&C9�ی!�Q�H�6�)�HJ�KA�ʨ�BB��D���vt�Nvj�c�܅�����]�O�?U��)�X6�;����fTC���A��L��p��lŌ[���>�)��RS���d���Cu᝺:��fA�9jUJ7xD�k�,��w̵0s��J9���e��! ��#հ��i��D���aY���x5����8�nf�=������@z�]G �Ј��j5ܑgS���H��no��ɇ-�h��ׅ�)̟fN3���M���8"aj�L�E/���\sU�r�ԥ-y�����v��o��&�Y�Tz;�I���l.��)=Ǳ���9b`˦Sҭ�,�h��~g6�3�V����k��L�=@ӏ^�����{����w�>tf7�gN�yn���̀weٖ�m.���������A��}�^�^�80f���&U5���ݝ���p�c��ɠ��I�Fv!�:gH����»�\�jfͬ�+�՘TZ�x%�������n���gU	
��ZSz�|A��<�N�����fn�j�4t�����ЩP�7��c��9̘w-N�ճ�L��?���ʊO���|}~F͏��Cs{^�j�2�t����Pjd.�0e��G~>Z�S�dݼ'M!�zwe�~i�{z.����͜QJ3c�bp�Qhś��A �e����kmf��˯^i�Tu��oL�nbJ�w�X�^����nӃFZ1�*�:t�~l�n̹�d��W5;×a�nS�r!�c6W��1������fzjIv��v���׭,��婥�f�]��q1#9�Zǁ�]�UV&� '#0�MRʤkO�9�L�*B��͖�ג�����pv�t�]T��rͳ��f�ݻ������Y2�k^�r�һ)y�B�YÂ*yoS;�{�p�����ҙ��u9)ο(�Ac��=K�-�*���w2{�۸�{���2(�w�����ه8��;��7y�O:C�/`�ϋ��uY���3�c��靚��2wb��r�5Ý.�;OF*���9�V�.��w�S���1r��13�Դ�ky��+����gk	*���v�4�;�h�Fi�^�;��.�t�ۓ��ǫol����%Y��a�����`���۸4Ѱ��u�Y����L��b׶'f3��o�p�'m��	�v�"��S�b�+tC�;y���5n�!���"ہ��5i��
%�عf�'���i��L�&R��AH!�IRP!Ҥ,�`B-��&d��1<�5n�&�S9tTc˸���H�[�����(*�d&܋o4*Ń�,�H�(�L��Y-Ƣ��$�����ş��D��tj�F�;�z���OfR�,�O>���jŸgL����9%ģ�
�+�P���x��K:���y����;�F�1�]G��C������{׮^��骾n�/2S���wGG2(�8Ԥ���K����
��ʝ�C�,}����O�Nλk���c�uv�7�ff }:Y�4��+&�|ݜU��&��6R^:'R2�s��$��*��o!�8f�=v�Խ'6G`���˛N]j��{t`̽��԰��4�a����S��w��K��\�L����JG�������5]�ݶ�Wrٷ75�s���~5����{KF0���t�	ğ^'���I� �n�ܻ+���q5n�:tnvӪ>����NX.�=�{R=�;�C��Å�d}7{����Zb{��t�ԚNd�TY�7��/h��ïf �u�{�س(?!�9L��־U���Ϟ�`@��tD�tن�Cg�b<����V����k���TQg=:5.�9P�צ�1�0��Fݨ�~W����S�B�i�M�Vw[�A�53�$�7�K���G��Y��P�<�^�֒����@��3gB��;vHn=w,L,�W2�LG�ш���T���B�X|�C� ���Gq|��5;��ڻ.����d�.�Ĝ.��Ʒ�h�ۼ�R�͌,�1tًQ��V��w	h��D�)�t�@�8�%�T�2��M��AM��m*&^�2M8�Z���"a��K4���?�O�	���(]H4�)spцqct֗ �ne6	K,b�m��ėR�y������fm6�**��.f�Y2˱��c]�i3��I@�a�M�����ʓ�h��ڮuɁx9r�Vd-�
f�K����ʸKk5�0�T��\��
ėb�<m��E�p�m2@W`�����~��[��[ųEs�ub��ם�%Ŷ��Ð��M��\�ЃR6�6�K�0��.�f���д"�����Q\尸bV$Q���lB�:ֳ6SsXL�/�.5Z��n0�ڥ "b�a�2�˭r�/ Ų-��Xb�L�Q�F\��b��L⃖�Z0M0f�]�ET�:-��� GA֛��U̱�ۦ�UcW�b�΍���� 7k^�&{X�4�Lюyv-�\giv�3�p��ƨH�ŗ,k����%�i����6�QФG�W]���h�����&n�λ)6�,aFʴҫ6˜r-��s����KY��cDy����)�nL-�˱jإ��Z��CK(����5D����8w8-�ljbb����RS2�:�P�VY���Z�%v�m$�$m?#��]�hL3GgeJ�
v��f��.o%֚�M/,�T� ���S-*�P��Y��3���]M+H�4L�u���iTؖ�fQn�i��Rl��% ��]M�f�-�F�-A�K�BMj&�b;k��k��yk4\D�Ѵ����!S@��^մ����U�WUZܤV���k�mP1�P�i���e�U�����֛L��Sb&��)�P֗�,l(UJm��U%n@Ů�iJ�CK���90�]`ѯ4&҇..,p�`͗�Ō����-Ι��Ң�L(X7�4��j�֒�1��r�#\-v6,�ݝKJh��(��J�mt:7-YRk�R9n�^3���WRS0]�d���8U��`�v�L�k�ƶ2[@�ٲ)vU]\ �G[t���d�b��
�ŖK�Ci��Ӏ���,�6�(f�]�@�u�gCbDE�n����C��icvU�lĐ��skPL�uk�iu�"F�np��z���n.�l��h�e�eL��8��$���+S7Ni����G5�+u��q��k�.6�l�,���Щ��.����6�A�1�.b�� ��tM�hYmò.�V�ؘ�u#4�2vqkkH�u�,l`ninEJ4���1tFf۲�����6׊i�
ͣ����(�bBrb�XY��a�]�;ћCC�Rd�Xư�c6��H�R���+�BZx�]� -�LMy��3�AD�Ph4�Y[6#Y�v�an�E�6�L��f���.&-KcV5��)8�ce��hɳ�y��`��`Nif�\��܆�GE�X$  K�QK;��fd �������6f�7���%j�K(����!H�1�1���6 �o4�h�\�6��6�:��b�^$�H�B��0Ȍ\3�сr30f�Vº�%i�f�H)��3�[5��,v��ʶf�jR��*`�kun�-���c�?7�xv�B>�}C�ʔBB ��_ �	�^�U��ii!b��H$�I�y���,��Bi��**��I!�!�+	1 )� m�,$+�qP��Hii �?9�3l8��q$%a0!Y���l
���!8ɻH�b�V�&09ݘ��LC���m6��BbM��e@9l�@<Cn�6��c'�4�1I\d�M��� x��yd�E�	եLI�m��1Y<�f���8�� k(i b���6�:J��gL�ݝ3L��x�d��T�X�|I�	�=��P6�o�r��4�:@6��4�[�5n���aY<d^0�s,��N0�/i�6�c�FШ.%{坲]ގ\@ߛ�giӜ�����m��k2��G/l�6�I�X�a�Xi6ָ�w�8�o���;���\��Ld�f��3\�/W�:CN��ެ�e��u��y��)��%}D}e�m1Qq�Z�l�B�/W[�q�:�����MK=�^���g;H!y���x
�xLt�ڝ]j�3�����u�t���g7kw�!��C���9[�7���g��'}^�+]�b��M� 3D�(�a��Ψs��'u��MC!ʐ>I,�E3�_ne���4Of�7�;N����wsu�DN	>R�a�sN�^K����G�`a���1-��E��-S
�&f����sS4�~�'Sp�j�g-�F�����7��D�q����7�-�$�d��V���(���a�3t+��'�vLZ�&�0����(B��#�N� x�K%g�K��Ȁ���l�g�(4-e����f��0�'K���[�U��#�����*5���90�}�Ϟ��'��ӯ
����x�)ɳ>�ǨA��C+�}��ӹ�Ć��7ro�DiF�G�BW�ͤ��z�<d2& �XC�'�K�o��j��+��{Bn��>9�������*�̢���geR�oū�9`ĊR3�q�����{�)�����ʡ;�7<�S���tZ��;�h�"S� I$�i�_EVjLjNgg/��{6	x��hʩ�pε�PiÐ�:�؊%&�B4�U�#�i�f��7�jɳ��B�92h�4?�z6i���V6,P8;61p�h�ie��Y�:&q��d��3p�+�ȇCsP-��H��0u����V%i�������ʪ}��]Ej�cc5�֬,�d$RŋRL)���4��nI��5Ԡ�	g�8C����3�)�s�QF� �ը�~+�fn��W�{qoX酄���@���s�Ϛz��ѐ`I9x?$�G��6d�
���U�39�M=L3�B��$�LbR��P�|� �2ӄ�n0�Ã�̅;	:�P�XHxº���c���аn!���=�2+�X?p�Ŏ}��ӧH0�6��U�u#����¿W<�^�6xn�kq=�)=�rRi��YXJ����:��^��f��	�b�2��5�[lŠ�GCLs��3,�v��YC"\�Z�JX�s�HE�Ĉ�[H"&l�r��X�Ƹ�9�&�.!sE3l��l�`8�X�di+��!)D�;�cTڜ貛B�v���Z�Eq��!��gh�7���/2`ґR1�m-Kr���"�#hut�,�lk	��Qr�Ғ�c�F�#���e.��Ά&�. Li�ãe�+�!Mֶ��4fhD��hg3Z8�157#�U����)n�c4Xf�dւ(�����K��6PKYIH�3r�K-��p6��8��G3m�'9'';���`��
H4�$���B!*I*�%HTY$U�"���QHd��H�XA@�(1�%B�*��I�'O��Y<�/���&�5�yĸ�Y�'$M�L��$�k(ieT����������=l��f,ՅF�kn�N����ee��
�:'����?(��	��:@Fu~��(�������r�z�5&1>8��5�hC�l�.SL�01D������8����<d�_����Y���`�Q"ǅ�B�[*�b�:����aXW�.4�CeېF*�{מ[{0�h��*�g{�{�:T�E��Tv6�!��X`�IĬ��Y5�pHci�Nzyx�ɨ>��H���0�f��,{<�|�Ω��ѕ�E���;-P�=Mӳ˗t[�E�P�j�î�O=��7BN �[���X�X�݁�ΰǅ���Ğ0��a�ՓN<�u�3�ǌ����?W	8ggϮS�E�'\�&��ŝ�y�f"�>���`�=�n'���Л�c��=μ�s��^�8���D��gH��� V�XV��y��˻��3FC}�f�C��v�k7����*��=�h����ӟ��?�P�զ#M�S��C���:ʋ��1�7�O+a��������}I�6I���������637�$b������{dǵ�R��������
���^���{��o�4�җba����7A]G$�0��P$ri�d�[��bw��ȥ�I�N�igW|;����,���#�$B�gii�"Hi���z��]r�0d�0Cz>{a�����Ĩ�D `?"�74bԱk��i�4~��@��^�|�;:�-s���2�����8}I���I�!�Ⱦ�f�RR 5�C�:�������""���6�F1���k2�;�w{�Y����u�Q�j��p�,�w�.Q0D�L��?
k�
�������t�gB1z���WE,��.U9�{%k}E��!Ұ����yD�r��A"H���0Ok ����t�sb;�C
��w�Z}��R����t6��b�c�z��+/cY�EYDzӬ�Q�2�dʶ�b~�t����H���1 �ۀq��,�� �z�� 9��m1���0�^�تt7��\�F�n��D#�hZ�i� Qi@뙠�a,7H�9�1��,�3G*� �d+_._!�C���)$��C�s�� ���i7 ~�`���x�2�q÷%�4B{��d���y��>c1�/���������	K���:YPt��㩦�
��A��"�rXZY��R�m2$��a���F;S0t36��Cm�&xʍ�W8
I<�:	��*$4B
#���Ԓw�	8�qu� ��GB�'�_)�$@���">�~�.��$:�Z7I�2��f<���N��P5ˁo�d���T`�J�YE��EȞk0<��6�ON�����p+HV����f_�A�H���˯�Xٮ�|��c�Q�f�.*�<��%���{}^6�i�A2�J-bE,�~�zm�6܉^ҠVa������h��lg״uq����ٿY。X#1��0� 4X����ɢI�p#AB@�Hg;RO�hc� �G3��T@�:�r�A�ʰ�8�Ġ*'`�!si�BIc��_},�����P
d�p�f�?K:��E$���(l��K��Xμ��FGN��ŷ�d�O���0�����$�0$�6�X��т�P�:t�#wY�,4�$�A�E$냱!�H/�sow6ޥ)�z�[w�T��i�}��zq�4�&&���i�6&H�;F��h��8�ȡb!D�)�ܫ�P��ipȝM6&�'m�8@�ET���VB	a{�����]|�ߓژ\�5.�ttnku�,>�~K�Q�=��#��a�9�p|c��}Y�R/�0#ӆ>�a�H�ZĆB̓�G94�TN��H肋M%Z�����b�4��j��$П��A�%S����"�E�;���Mm��Vf>=o)k3He�Nps`>�	7b�H@��8�5;������kbG�׿�(�Ts3��+���ǃ�0'����A8.�G-�~�F@�wkN�p�� e�M�����@�V����53'[I� �� �g���S�ՠ��!(f��Â�3s�ڠo�H�� I`ΡqU�(�;kM��fB�������c�8��:��	IC�<:c9�3��,����Z"/�[��kb!�*>��l�5йf֡�����9Xr�� �Y�7!3cIk�#���Rܶ�ZUԔ6�vn93t�J2즎�l8��/���s4
BJdhB�~�������S�b���{��F��Ү�!I@���0�ub>c 3xu��~�IP�L�4�O!@h��� �|����Aǚ�l:����F���p����rF>�Z�lBEF��B�B�D�6D���9!�'zoB���F��u����<���=�uz�9y��Cj�B ���4�¡��~�̬~8}�{v=�R��:���:W�x0hv��	@U4)w7��1,o�%��P��"d�X�9	x�!E�I���1r��L �#[�Eg;i2��	0���	�BQ&EF����i�E �������6��z���JU9�����UU�?�7*v�4��l��v��vQY������D鞂F�SI�2%C����?�@�1�?�rt��j�7P�~9y1,��0�����[��\�v����3ð�p΍��[�\dF-����
��]'Yy[���{��(�R≁���6�_w�g1-�55{X��)`5�zA�UNMҵC��t�Bw[�&(���eIt��鎙����񬠢['�wIoĒh�ޮ���m	k�|_%.O��3i���{}���x��>���j�ٷډ{��%�0.N�.hH�{��Գ[yw�J�NQ3i,İ����B[���E�H��I�1��R
 �,QE�"
� ��AAAV"(")(�P��)b�
���Y����0C9�L9�κ��b;�� ��Ӽ�t$}����$O����S��m6�p@�>�X���G�]LaS�KrA��"æ ����!�+/8�;��/JTX��0L��CE�vP���$�	��׹��/�1ƺ)�*�=�֭u]���(z���D�)�P�/�yB|���ޏ�d�fQ�Gϛ���l8$S��x'~�x|zC�5�,�V�&t���b��Xy��Wf$�oᠼ��Ģif��a���ް����D��8�#PB:��O�a~�� �C�A#��>j���&�z����7��/�W�qe8λ����e���#�HO�P�D�k�[o��i��*�``�c���>�]t8�@:���Q�<�؜@��w���E�\�T���J.ʤ�Kg'��Lw�,!�>�@$A~�'�;�*E43����.fa�p��*h��~za;�����G�'���S^R�ě9��_7��˲��N��� D9���D�+��4$2;���>��n�@:��0,�R��_���ڋr,�#�`����og@���dJ@dac��4���A���[���{�t>A ��5�M9C�����!@�DV š#��T#��l	 �bT<;��)v%
�!���{�=���eZ��"�Gg5*�C�˓36[V�S1eF06� ��	aѭh
훶m��0�&E�V6�jkHh�&YL^e-�sr^Tt�8��'9��Q6���T��(���s�BKe�I��N�؆&p��I��#�0��Ms淳�S�<��Ja��;��zv���bT��� t m'���!�T���P׮�N�Q���.R9����A �o��ο����~�ې-��/�E�����@-��T�v7�p�q���@���kb��Np�l*Р�ك�"ŉ��K8uƗ2���`�����zo�������P�찅��zQHh��2~���/[f�6�����V״|>�k���0�AY��XX,v��,�oE:Û���ǠW�{�hhУ�š%
��/�f� kؒcQ!��*y��
�87D
���thΐ���9P���.0��p����r�ϛ�$�>�}�9�3�u,�{���X�I���b��!Cz�������A�ӳa�=~������s���/��Bh�q^�)�h�2�Dӹ%Q������H>A�q'�^%E�w���QPZ.��w���3��E䞶Ӟ`ގ���w��4VXT\�t�Yw�G���G�Hb>."S	���)�0�O8w��R VH�a�0Xa�A���T�dP��Xv�W���Ƞ��&w���|�`m�P֬e[�[�>��v P4=��6�RΓ��aA�Q�ܬ�_���a��FG�V-�v����G�H��$��ԓ�P4']H �	��(P�gO�kc��ն��n�f{��~ ;R�_Q�X7�p$x1�O�`��.�A6"�G�̰�cɉ:�1b���M	Y�d�(����p2$L�i�T2�`�ų�Sbtf
�ֈ+�	�c�B��'��cE�sXPX�0D�r9}�;O�3�T���bre�#���߮��{���-�"�ŉ�i��W�l&ı�ɦ*iu\��ݴX�Qҍ��c.%Q�i�Q��,4qx�|�s������:i��W ��<*�=Рp_va! �g�F�g�Ҋ��F1��/B�1����T��������C�6�ë���/2>����"gu���&=^��@2�.�ЁFI��P���$EФ���,]��?�(e������͏4�a�Wp��2��W �?^��}O�a��w���/��#N<wm���Ę��#����*�'bT��y{��x7�X���Uw�i�~ =� !�^v *�3��7����� 0���X��Gm��!�zn����T�&�h�����!EX�,�<����-49�aC���w1dT��J��Ӱwc<�mC1Q�@]�@Et�-���}��t�N���P}����dz�	�Y�
����Q��a����i��a����m𿝂�\��9�LhW��b�^+YF�\�!q[#eΚ�������xH��QB�^�!%Ǭo����uc{�A1	%�>����[p��j�1�u<;��'߶���0�H�K��m���>#���T�v���?f�AԂ3�}+�M+�����aRn���2�$,L���j]�(p]�=���l-��D,V���8@U@��2u�K��
V���'�������G���9�&(�e�($+yqEE	\䈎4!x��J����i�CE&�ݵ�4��]�|��-ł��N8< p�S�V�l�������x�B�&7�(u�ձ�x�E�ϣ���������y�7���KdG���
�]`0��_��X���H�˱�1~�q-��o�X>u�Ű,<�̌��u*��]׵�_d�����̊����Ʌm�ݑ�����i�"Y�%@z6sQiՙ-\��>�]y�ϖd��S��j�S9[U18KX�����uQMNVl#�F���ߋ��sS��[�I0p�k[噔�g���S�7������x�d�*)�R��p`�6�!nJ6R�t0�DɆ��sTѵ5�!���moҁ9��&T�+#(��OA����K�>��nOnk���&�8���q�����{��	�Ͽ>��6�	��X[L�W�i\,���SL<Hj�Iiae��WUa���X��R30Jdu]��`E��Fƥ�:۝�jlMԪɍ	un��\0宎Ԅ��?H�q7�`�e��ō�Z��^�����s���r�2ؘ&k�"6G����lvb�QhMH��i��٥L�T�e9�6��T�Ä@�ѷKJ��SkՔ�LУnHDٯ
P˱�ʏ	�9p�2�mWR�ٵ�7�X[.lf�;��N�f�+�&��%'qkB��:�Ab��Z��e���h]˄qs��a1s�T5+i[i���.��*�s��D��$D"�P �I����A`,R"$H��U���
�E"���X(�DdUP�Y�ﮌ5\�X��]f��s.��Dj��kA�7&�pj.�ғ&�CYu2�]�]3�� T�l�@�#u�&�ӮH�ttZ���.�� ��"m6�~|�ƁC�D'�PS��8�a7Y�`�"���ޱC���� �t�9A��m�ւآ*1��\`������h�^xdAm���a�kF���(zX궙�ghؖ(E�h+�F��kx~������[�*��5�sp �Xz�}����=��	�HT����0�:�	���c�fϪ�L�*��p�e�'���[��XC���a���3_������S�,6=<o���,e �J��^}ÐN���(��<NG���Ly�Ш������N°��i�\'�j}�MF���Ц�Aq�ǧk$HѿY�	RA	H�x�b,x�4܉qB�{v�ْ0{�X)�� ĥ�Q����t�������a�����	�iår�NkE���؏@��)��Xu��/P7�u�,M�ǹ�!sf��р��@�a�r,X�5ȡ�:GD?�-��B�Gi��mٟs�����xc���3/�q1��7�Kd���((y1#pa9�����M>83�A���m�F�ʡ�B߰AX.7:�M��8�X��ZE�R$G��^(���0�>�[�ŗBX�-�=s���2�6�O����:={�Mf��c���������/]�l`��&BE�j�x{�#�E��X�Rd�ޞ��H�N�vM�
��3~|�R�8p�m������m����Cn��0X�R���貂�AǍ舑8F����s�Ц;;̦Ď82p-�c=����M��[��3Y/��oQ:���brb�;�s���O:xr2�E
�����v�*�lG5�lK�4�-4�.a,ɢ�e���Eq�aB43e�12�v�ϋ�S�R��:����T��(ǰs�)=cjh_��zr]��pzf���K�E���FСP(��u.�P���8!�m ׎I<�{䆅Q�Ͷ�6s����x���F��!~7w̷g�)b��b��hu�{���w6sH�]n�LW���z��TdT_,#b<^N{o
O�+��ֻ��UV�b�w�F%��&����cd�.~^�$,`�&�Pf4r�T7�-��&��P�wP=��u@�p?���F��]�1-!�jdXBLq��%`���y6�d�=���X�"�`��j���z>�|��%���&ƃ��\����T}<��I&�^/Ƴ���56��<�k~;�_�M����t�8A���������مWFnw�X5��RfΣ�j{!v;Fh�R;�AT���^-487��^>�����>ecH����y��O�[��1���apL���a
䐑�}�DFO��Щ1;��Tk�N�n����R���-`�+�b�Bz�sI�#���h��*�b������ߑ?�Gߗ����zC�71��֦�g�7(���22�+FW�|���w߳�~��+���-����t0;�E��*��"���}���TRI͌���g��?_ڷPtE���]ȧ���s�
��8*"���iI����p{�/<�Ae����<Nq��b�oh���μ�\���zX_)W��ل%M�0#u�qeQ���_4�k��3UZ��X�F킁�0FҸX�e�ycm�
W��gmX(�l(Y� f�5� ��!�W�á��ɵ�l�4X��ϱ�r���cO�K!p:$��m���X"�Ur=V�����R�dq��s�.�q	�b�n��KH��� �v(*�7#o�V�'Yl��h>��PL�V��C�����g
��(��#6T&�$�xpb7�hr���\��B
!��%�O!C���S�S��xfj��qR ��R�� �8$�G�����P���lI�B��c/�;�#��fdfT�M�a[���n���������m����~��`�9��B��%l�gF#�q2ҟ��ˀ�b	�m����~M��'LC���`��o���u���l_b7#�"FH�\��_����^����|����B\�'Rbj��ID�f���ݛ�-���F�Q��[wn
iB��p��;Ԕ�����̙�p�n��m�םj��޺'_�G�o����Mm��6�˘<j;��{�;�B��cH5�ų�"6�m7:���([�lM+_99M\lY9y+~l�k��:8�ﭓ~��!3�CI�����Y��ٳ�;���/ݽmԎ�Od&:j쇷�(y�{��4(�|�9��F���$�&x~,��TX�"�E�E��A@P �U ����R,�$ ��2,#����~E?�
C���aU��B�S;��3w|�x&�Y���;Ϫ�h}dUȘ�J����XiA�(qat�eY���|���g����^8��f�y��6�.Ǖ�"C	�d\ym
�z�l(���xPp��>1?X�p�j+E�����([�A!�_m~�x�����{Odm�,��?N���6��6�b�\����Y��;0Q���|!п��m��Be&XP<=VbǇl��Б��=y�F���bb�+�Dzof�W"�j$XB���#n[����,r�6���5c�=�1���G{�X1ꩣ�;�4^@��1.�{��>ڱ(���~~��P�/\�9�a���w�\��.h����;�r����v��%i]FWMnuj����a�u��5�r�6�ƫTeu׌.�4x�Mp��ЖS3LYvԕ�3v�k0����'�������Yun��&�';³j_�Du�c�'�tBo1��E���#�C��r�ٕb�Y�z�y���X���
ѭ�ԯ�m'�XCgP�^�Ѻ�z..¾2o��&"Ph�TC-& ���wd���Q$Hj�{�W���pE<Y�ӟ�F`5tʻ�xUС;Y�b��3~�t�t]���po��^\��Ep82<:�m��=��N}Ϟ
�U���mh�[<]`C)��"�s�b0p�5:�vh�	"�Ȋ�t��Ol��/ׯO��s�g6iF�a�`�,����
A�Ы���M�+|��O{(��z7Ky�,!Tfv��6���#�R1�
�(a�����,d;K2LbY�n���ؿt�A�{��Bl��v��	~�`��C6z셳�/��-4ؒ"����btQ�,���'���+�#�[,af��0�m�����g���a��Y�����5I�B�3�\]X�\X�	�R4Hۚ�i9�bâ�["�|��|ű^��S�������ϭO��=¸#��&���L��g)��Sw5~ϸ��{m'�sk���w_<�����C�|>�b&��m3��cUħc��@�3��Q�ow����U��I�ܲ&�w�)����l
'��6\M���S#�C�zl��PO�رn�m9m��U��5N.!�h�b�e���&����6�\`���*k���O�\��nЅ�C�ܩ�+oA�e:���LC	(f3���k�B rmf�����еnњ���4*�r0�mt�������e��(aکUn�ZU2�R��x��x�x�{��σ�f�<�l,v8H���иV�bl3Q�̰�`���7~��ဋ��K{x���ƅnȐ�u(�}�A���Z!��t<�xx��i�o�3�@n�0�Wh���	�#�z�����(p��q�8���X�bs�`�}�a��)� �L]��lf�;�(	 _�0s���s(e�`{�6�v1�cB��&ǰ�uO
	X�]xE�[���ӎ�Æ��J�Q��&*�o��^}��]�<�{��7~?O($:�V�[�Ga�0[i=�J�$"�:2zb]M?rEKm'bx��#}x gq�Bhh����s�O�Y� ���@������U�~��9��$��-θ�f�𪞟@���z�4�4��̑�%�09�b�DM�U5�6D���i6)P���s�hyn	W|��'Px�(�!��M���qM3"Y~*����y{��:�}�COퟰ8���B�=���OxX�<`�����C�9Ed	&�����4бUS��o��LȚ��&ג^`z�m襆����G"�a���ykLx:u��N���	��
}������}E���u�1qc�u�Cb<ǂ� �]Cs2M�+�${q���D��>���3$�{]4��=,N� z�������ǓN�v��^��T��RF��7��{�ƚE���A��d�Co� P].w��������?ܿ���{��"�ӟ-N%�S�mv:�qN��Z;4Û�V�r�!����u�M-��9;(�z�(�ѣ���<=y]k��V����g��s�Wإ��v��&��M�7wnV���N�b	z�F/K�n{}�I��m��q)Y���f�|���U��$��ç��T����^Nmf�'��(�3T*Ŝ��T��+i��N�Vה6nNA�y�x��s�|5oG�r�����޷cv�ǻ����{�ٱ�VF�[h�Ђg�2Y���ř��^b�#vƸXG���v��\ڐ�'W@�R�͌���8�Z!]�B��	M-�C�E2�vKl&.�՗%���V�SY�	K1�	bd�;  v۳����k)/l�#
bjK(�cb[����dfE���xfmq�#U����AD�c�=�a���űlے��j(S�l����+��M,`[V�[t@D5�T)l�]x�h��XJJ���q�H�bܓd��pm,b53�XYj��	�l����a�!�g^%a�)-o.dE�M�W;%�"B8R�]�M�&�YG3�a2���\����AHAA`��c �()$R"IU��$	N_<�]s��y���\��DQ��[@u�j����nB٦�nv�`w/-�y�����Y����ۓ̬W�:�Q���?U@���-��V&~��|�{c�[� p����cjƊ��Ē��hd=�7��/�����"9�����|'��g�gw��ɏ1r�W�S#Fv���~a��dh��@��k�A�6��e�t6Qө����:�ǣ�sô�	���S�)���؟x_=���i���7e`ٕ���0��S;&ā��ϼ�BDu��z��\3B��+��& "�Яzg���3�:}B��Z��B�C>
`G��o�{�E	&���ϯg����q�R�Kn*��X��MlZ��{ٳ��!v`(�uU�"�V?P;�,����6ت�`�����M?�"a���/�'�ު�y>?uH�\�6��P��3�~�7�x�x;��UO�~6��||;���~�{��_��-
e��b��S����g�*���J�A�}Bkm�l���k��49�����~�G������,dP���n����e���ɣCW�W���k��:1�1��_t��K �m|[�����)?��pL�݂0{�b�o=>Teu5�a�Cf��Ũ�]:���t���g��3y��\�^i�%k�S�ۧƾT��;�
f�vy��_B�t`r��`��l`�|n��>P��T�%��u�3���m�
yX�z6�Ǌ�pd��P���e�{ð�|躬ۣ�#�A�혡�A�%]�%<8���0��f�XV��\;[�喙"F�Ye4��a��F莨F�!����ΦՄ��`�.D�z��m�ĸֱ5xiuΐ�(l&Б�9�/�X��U�}�aĈ��<M�!TR���ЫP3zmf�X����B߰N���;j����`��n�`��CҡP�m�-�B�h�pU�s�w03|Q��6�l��K�2�:e�ʾ�k>w���C8@���څ`֡���E���9]��z�*�%ŸI�̪F%�UF�r�_xz(o?]�*�:���n3	l�+$@B��P��bЩ/RO�u���b���EtP����4E>tRz#~��`��"̌(�y���a����d4�pM��3ߟ4��;����P��*c�b�Z�o��Y8p�wCA�N���BD
;��߃*{k�~��T�I=�T.������H<{���D�m��AR������{w�4[ā4��;xC%{B�b��SΏ���������&�8q��+֎Ph\2�fb��m�U���{ڒ���dE���7�b�����Ym�ó�z�_M�ɡ��Sxq��x���މ�?���f)'\�MMW�Tꦷ��t��p�b���#����	`����-�y!Ci��=]��S*�Fwz� �����4��걊{60��oG�X�{K������&��M��j�E���GhC�lz�.��@����I�׻ϊՃ_�����6���
ʏ\���n?6�'�9���`��pH)�Gzhˬ�\J�d�;Ȓ�?���~O��l���� ��6h���l ��i���"9�`�]�Հ^�i[��pf+ �F�V4����t ��Wk�h]v�(����w�%&�{�F�0T]��xŒ�ٔ���3�Hx�D�%G?zpZ3����IU���P�rk����^:"+,n��m�h���V��ƈ�^}tlw�&e,eБ�������d��u�νr}]ڸ-5ˮ6ʩl���4T�ed
X�Y�8(Dh7�~�J���"�'�j�����a;F}�B=�"ì�������[|P~aH��'�.��>h�$v$.}�HJć��g�V,�c.�Ў�F�4V�������p���&���K�Q��[ne*�J9����{��{/X���DPr&���m��F��̭��� b�=z�r'�~"G����?|�?BW�/x�O�?үc)�}c,k�Z�����\���j���9u����+�b�=�p���ǥ��b�qL�T��p=z$h�0e�v>��$d�Rf\�<	^������m���o�U��Z�s�t�؝�)��J�T��Ŵ3�ܽ�]<\��{5�����;��ӽ�xj�-�*�mm���wR�g^�{��zƵ��7 �0�w(�6�k����Y�e�`��t\��r���3]�E�g/3f��s~�� ��" ��"�"�Q@U�*�Y@R,"�0�
(G����3�LԢ�P�x\���OW
�u���xd�{l��X+��I:љ����A.�}»�	bD�	+w�G2B���N��76b�$����0��Q�=��B�{t��?��5����x�r(/����!-�*�Ro���K��V��
#O`���ȏv��Eb�������:�}��5�{�f���l;�����Tn����sM��^���`#��
�w�w~�/���L�e̳-`&2�Sc�Exr��hg�b�LV��|��b�3S��n0��W��"�v3�dH��^|��y��.{~�
�S`�zx��ћ<6D�c���r�3U�9�^��T̥~���9��É�6�����;Ϲ�Z\햍Um;5�vN	��f�*�)�$�F�r�<G���T1(1���)��c�)���,���.��]vn.����~X<�p"e�d\�m�:��m��3c9�c&¡(�S�P�>�-�.�
�x`��#���T��sžYb���ؠ���t�+M�`U�P�w��6|��|�O;���x���Q�-�����Cmد��9dXǢ�|��z=�\��d��sP=��M<�����H��[�kv^���.2�äY�W}� ���cm��������PC����I�Q��p�^�b�Bz�sF^���S�~��4@�ŝ����1�ƞO9M�ͦ �8�.�Y���~�ÉI�FDP�;�����}���厰��nǅ�����B+�s!9�^i6,`�xO{pGr'ι��H�S�3�Ҳm�٭��wL�����ޫ�8���G�M@�X˰��0�����k-���r�=�%�!�͎��<�~�q��]4Y��.pe��x�ϐ�>i���g������OO2��v�0:�M��u&n���m�8�`�Xĉ����!#@�y"c5��<���w��(Z����3-@s#�:���	�%CwX-�[��u�܊������:'^�|�}����y<�~L�c��V,r+v��G�h��"�\1���*V49�c%�A���� h��bE�8/>����T�Q�aUG�P�'���)<g0z�`�`Ov5)��M�c�g����'��24Nb{��,#�����9�i�08R��[%���<X�,X�i�2��,f��k �r,�&�i��5�p5��m�tݴ[���b��*ɠ�Ů,^���9��MMvI���a�x�vt�2����2߇��v���Gl{���7<)���E�p�r�DH5���P�X�G+�-;L�+.��BG�o��0v��&����^��bfdO���#���\4��:�m�A��~��=}��o�M^s	4,Z�]x Fk���LH��yL���Jw0�I�Ѵ#�",0Z� ��s�t&0+��ק،�ca/�bD��~hp����C�x�W�8{m��X���	I�Bkފ�ϯ���!�!�K(�ι�l����h�l��^D�����E����{�`ߦ>.�_�F8i:�
���7����t?�d��0{pU�K�Ff�\<
�����x�ߠUja�/�`���8)�m7`��١�:"����<�z�ν�|����].�����&�Bl�����;֐�t"E*�N�Mн+wEE�l@����:�2�D�ʳr8<��:�gy��*�z K�|(Ե��)gj5��MF_�iLґ�	^S��&#�U���E��2=֛bn�7^��|�_w������]Zapl�Xa3���'�����>�0;��Sbǖ!Ǵ�� ���l���b�Uq��`�LW�N�9�vE
��PΒ�C/;����p:�ޮ���6�0xPl]�_@�����>��+ߛE��~�+<��w72. ��#�5�5j���QV�Ǎ��������k|*�c]���L9�M.Ţ��ou2�~]���K�=���Z���ƞ	����w�|]ܭ�Q�춄�n�O<��d�<�y�e�c�2)�%�{%9��Q��M�W�^m�����Ӷd`�og��GK���ބ����IbE�Ͻ�o���|�ӌ�Ҹ'�:NC^W�1��k�{����v�uX;|嚻��t����q0~E��ZiQ�4�R��r1�`˲���)Q�q���i�a���#b6̨'X��SbeR�6]˝a��]��ri���n��h���jq������6�L����C\Χ3��%�"�ޫ2�ڗ&��lhlA]ck���E�),X�T�.�9�
/V���aH�ԗ[%X�k�n�HB�g �6I�U�Il�%6�����F�K]
�+6h�K�kuZS-�Z�B��Ѝk��,1\i`L�dl.6p!M��if��N�/l����Ev�ږ�l��++0�
��Jg��t��؈fk��sR�$.(�=H p�Y��,��b����%�Y�g�:|��k��M�1-P΂�a�5�f��q0D,fB��p��s�6θ6�К�#-@6���vF�B�L��b�+,�[R�pʢs��~z߆��I
ă'��)��7�!��L��^	��腘�"e���8Gh"B
O(�\X`C�^bI�0�[�2`����W�Q�O�OGo0ơt|}�1�nsR~�D2�F ��(�E�$�n�pr��`�{l�¼���W|�r03�S�A'.'�*��7w�=������$B&Ǉ�A��BD��F�3x�L�=e1Z�P�� eq��M���5j�t�c��Ow�u�̀[ ��#�^���c��D��^�'�ĉ� fk(��3��=}P��셷��,y�4��	����8N�,�@��G�Ex`��=r�<���½�ɉ`#�k�-�vU'������J�ewc-��2�<�Q�$`�f�#y�hЅ�A�Z���&
t�!����d#%d8l$�KpKp`��6�,�����&D�z�������SM��"�w{�#ك�����غm�=�'���xd����������ՏFo��B�o��)vcD�q�
tRP��S���F�nrO���i�;X��Ǿ�&luR��__����s݆a��ŕibs��VF�=R*���n�'�b�|�5��*���Ѕ��0b����B��޲ףGD���N��T�MfOG�E��n�m`�@��0"<T�7�����t.��������bvg�/��E&�z�9�{N�0�M1�\ƒ'18&y�k��:.��ud�E�3.�C<��6��VZ�]J���)5(ܻshV���5�b9�\m���qk�r���nD����v=����(a�i�6�Y�T���T���1���8X�j^v>�X�pѽo׾e6'G����)P>ξ������\4t��COh�K�@a�1|;2tW��P*b��a��b$��_����{��:"�d�pn�4u���_c:���s	�qނgùƶI�����lES��"����`s��i������hP�Lp���i�����<;�����c62��]���':;0bעX���C�{;y&`@��8	2BA4Zm�`���H7B����<%��華9����q`�'!W���	
���C�o�o�I��"�α�p���j%�¡ӓ/hl�`�1!��ހF��y��y[R�o�:�Ɔ
0M���u4R����H7Lg|�I�4=�m�}����SsCf5˜�ʋ��꺤.Dmz��C��Ƽdm�U�,L_�xHt;�s
E��eTȾ��|�����Ѿ������G��]\���p"���U�͎�,��}�p��ֵ2F�
�pz�H�'E�e�q1�ŷ7�|{�H'���ǌ<a0�l7�b`�[E$<���� �8����2���{C��T)�9!�2O�Sha �#��~��u(ǲ}���e�Bi�l�+c�m�
;}#+wA�W��&�v<;�?�� ���p�fK��6W3���M=�2,�IFV�ى��[��ڼ�C
���D[m#*7m�
�:"R�&��Mu��VWM��::��U��n��ӆ�͓"��Y0.-�B!����������-�,!�9u��l]\?�d����5�`��H*��v=a�'��(H��ߩ��w��Pw�l��n��3����촸NϑO�*��8��!�"|,g�,o�V5�S[+�'���B-C�ɅKm��g�^c��>2DP�ڞ�[m����f3+�6}5�l䪈U�<��6���P1�G����ۀ�D�2G��٨����lX=�^ثCjǽHbrQ����	�?wD���8�x~�>�����D�D�=�po/�A��Q�~��|D)�^,.7"�G�����2+�ˢ7����X���QR
�c{�b�SЊ�j��5n��U����2�A�͝��a�Ti�ΊP����	ˇIS+|��u��W/$�7�I�;e����G�o&�u�g%�����ƃGd��3۷���I��z���?{2���D���d��4��1zem�g�MăW
��wC�%�����om�g�d$B�
a+S����^��a'X�������]��)�]�<��7<��3�J��zb�����lż��^�����r�<���X�D$PY�Qg������lθ��Ē�>�DxOn�[ü��yEu)6F����:�����f��d�v���Y��l�����3���;�&}���B+'�|�qk>߻�	�B�j쮝��`@Cu׏�j���;��#L�����8G�m
O%����ǧ.b�/#�:�]����;�2���Yr|���d����χ}���P=��v����:�.����t��wц��]������z<KdD{G+�=p���B�'x�B�X�~X�볖bF���U��Cֽ������s�:{�,Wh���
D�烎lO|{A�1�������(y*B#(<��Ȣ�瑾�����3	]DK�*
\��ǜ%m�4�r�Ut��Ib�lp��-�nj(%���M��
;m�`�I�c]�u+6lz�L$�M���on��/�c��r*��^CW�5�x P{����1�e�8mB{Q�mv�
"U1�Ȯ�c�z�6oH2z&=c=�t-��|,lDDGf퍉�g�ZH� "�[��V�f������Φ�i�:�G�+m@�BxY(��_�]�����UbWK]D�ͪY!��3����N}^�X�����TgB��>��2Dv�q�a���z����L_Bmr�.):,O&�w��+E�!�.߾���[Ի\Vm�0(6������UL92y�O_w��d�������~�вD}^�Bwx6�U�ɷ!%��,m���9�l��+�P�Kڐj��NVS#8]�ʽ���Vֲ��S�="�o��c���M6߄�C�BBP7��#����l���+�����]n��hdo>O��xM<	Oc��f�6�`ظ��j��`����U������1Q�Q#��o�=��Z�%C=��v�윯-��u9=��B�'(�y�y��נuN��Y��	뻂�u�����z�I���nM6��,�{��~�ɺ�g���_���ܹ�����4=��w��3��y"qHN�l�M;��R�#�E��R=謥���f2�A��!X;��n��B���c��t�8.�_,�]�cX��Dm�߳��vq@��ߘ����F38K5��m7��E4�3�Ŭ3l7Mv�UR�����R�142g�֮f0)��4���G[�����u3Ul�65�￸o�5(��9�{�ٌ�
/��m�M����7�?N>�������N�},�b�J}a���'��\���E���=�=�x!V�n������)�P�(Tu^���	�迖��A�	U�Ճ���xH��|Gk|&�-C&��<!^�J� t	�o{T��1�O��c�0GV�:[��������j�phF��Y��. ȁuS˔l݊���c��Ӟ
���1�M0G���A���r�(�f�u0FQ��ȶ�������7"��=7R'�8��oze@P\DA�0\ʱ��R��|�u��'����7��#+4]��wy��_8�cMg�[c��WP���B�^���+2�_ٟ���׷�W�U/:^�{�p��{�(�+*G3R� �z<�{#��9t2w̷�#����5�+�o	� F��>Bl���$�%��&b%�<I5����&��??��ʔ0��?k���G�7�ת�x�фM���+��m7`�d�,����HP�d�ʢ��+D!ǆ�X�<G��Yy�F�Q�D��B���"̛bX��#���p,���!�nH�� C��C�=�8~��.Țd*͑kj��<�NLRK��X�������v]କ�=b�Ӏׅ���Bi�z��z��M{#�*�V�N �Ŧx_cR�#��o���W�c��"��n��ke��nm
�)�7���ڻ��m<�fvڬ����a��R:i��^�+v��ж[y�Ojf�/U�f�t�y-�K�|F�g���.���Oݱ$|_�k���g��xaP��)3�2v��ٜyFÔ�|4�M�����e_x2X���{&��
�3o4L�kU��lU���P�R�n�S���34�l��A�e���������q3tu5|�D��ٗ�,�Ϟ��C�pq�=�\LB�x9	��=}yߧu�~��9�^>�4��.P¥6���Vc6t5.]��mnm�j�\�7�Mu@�T�h`��&�^������4j���WL�j�\��PE\��͌�5�a]��i��hF]��1��4�s����g��%�X�GYYxL1 ;�,n�7ca��㩇e�f��&�5�Q���p�h$ջcGJ\r�͎J�����a��̔�69 ���V6m��)D�-b�h��T%��a�a�Z9�8�-�j�
��u�4�J"L5f\D��a5Hv��e�#T�K�\�h�,έ٧�݆�˦Ji��-0�A#V��M`c\��T��b!�-)���j��I�w��Y�n�\sF���d�դ�V��@�)t�'r!�3I�U�j�T�&`°�X��&Ϊ�4͘��i�&����#պU�d�	"�X��~ÆBད �#3ЊlUr_-�3�P7�>�,{�kj�M�ϨmU����~��(Sƛc].ჲ�mP���CB��b-�z�����������F�(;��8\�!B((���%KkG4�~cU��&+;����r4\h�z����F�Z��X�2{����]Rc��
w�H�Sr?6��˯Ɠ������H+o;�:��ј	�M$����#/���z�,���nE�Uik����X����!���ĳb��ZF��s�n	���M;'~�n�6�$P�AJH�x$7�b���V<Im��`������NytL�6�k72؏`�����,�ѻ_�<ى)�	-k�&���*���`���" F�Ԟ{�����lB�e��p�����	�Χ��N�}��CEC�k��|�@�����	d��C�0`��!֩m6�{�WB��G]p�<�q=�P��}ӕ/&T*�p��kso2��m4+d�w����:"~@�ȭQ�"8��}7(J0��P�m`u�`�h���:"H��u�!��pU�c;�Z5��
�C��Σ9ǚOD�{�� �v��cv~��W��o��bDAB=-���/C�=�ͷ��c"���BG �����yn������tg"�Zϕ��i�Ǉ+1�\�KX���j�JM����b�Dv%!��W+�6	�L� ����rS8!368���F�:V�d�X�q���E0'�k���@�o�Pۊm;�b�jo{ߊ�X�wϰW�i����=��!=�M��w�L��֠��n�k�#ۂ�9�;����M4&]�M�f�dm�E� ����/uX!���C�X�8��&�1��Ύb�~�?C�dP���^�G��L�uB��/Uw5�`d�a��G�\��qb�z1'q�)h����c/�!����m�*���e(>ڧ�C��&���7����x`7>�N���i�>�A����@���J�;�ih�B����"6�Wɧb+���b�t<�U��������L���X�õ��<�H�	G�}1���v�ps!^�=~	�U��اuc�|��p8Le�h�4huu�i:���
�>��b�}�z&�Y��߇���&Ek\�V\�6�OE�,F@$υB�N`�W�f�DЭ�"߁=�Δ������;L��o]f��y�$��ٺ<Eǌ�{�@��]	'�p8�'����oE�}�ę��v�7v%�[����׳׉6���y��?n�"Cqt��_����q��j�1��1��_s���x�dn�m��5o�-4.lg
�ݫ
�}A��ο4��LX�A�\�*ú@�rIl���|�B�q��G� c˾V8]�BCf��`�������N�ߜ׸ h�0��wpw�KQ����%�mv-t�����Z0�F�Kh2�\��W��Ĥ]�Jʁe�0s),qWH0������]�ZiA͋�D���&a6EF��C<"�z��ŰE��.Ĉ��f��y�@_���r#����`s.�"ݏq��� �s���c��X�����Ǎ��c���M縟%��_�]�E�s�Q�E��i�쁒/�7�q�N�,�����&+����q6�^�Vř�.�����5H���/C9�S`������V�(�Ȩ���^*���=�[N���VĄ�;��e��Ѿ���BGU��Z�쳂s�����	�,;%�I��#�nW2�p/�C��U��|jm�s��\Z)�hJu�'�1�";�,�	;M�|`-�A��:��ǵ���Ү�._�C�fܑ*~�ݝ;agG���_�������X����D�.���JS�k!NE};���qN��*���q2qL�m���ѽ�r�'h�09sLWf�8����l8w;�s}}K���C9ٍ^21�v�|c�����^a{�iĳb�\+�.�ɘ,�z�7Dh�]^`�+^��r�'�u�{6d���w�+��-��.�}����8���.����V_-~�����ѷ��]z�P�Day�����&���*;�P��j��9��4�^+�CW"b�O�hqCR<�c�ӂ�7Z��WL�Vu�i�������&}_�M69��{�i�"pHR�g�<��w�[dl���+������kfp�n,Z-hpu�B�����Q��eeH���뜨ɛ���\;<��������/�O�x��}��Y��Ba�@r�[���|x(�,H�^"kju��<C+iu[qX+(e��=�C$_��bZI��÷�ǅ
|&����i�bf.4�83��
f����CB�ZI��w@�C<7�;C���4W����jė헬��&�cUM��I:uRٓ$���+���w+���M�Z;[�Cb���iv:����s�w���D�u�M�����.�tw.���9�f5�r��p�n>$l��H� ��f��ڙi�hE��
�F�Kk��*�t��;E�!~K(W��Ya�/s�i�lbP9�e�ЪA�ަ7�h-7�w�P�ł�W�^�b"�}��e������T�e�y�|��'��)=w���({ua��\��|�z�j�Yڊ���6�p��!^/s�b�{l�����q���^2.k��X�?{�Ǥp�^c3F{ޫc�n�t:����~����l��,��C�T1IPL(a����A�Xa�Ϗ�D���=��x/�7�����ġ�~�Ք݇�{�Oy�����=:_������Y�®2��*�$_����OnF��s�g��ދ<P�>��C��i-��mՉ���xX�/�$8��G{�<�pR`��`DBN#�L�	��|�4��Q�=��Z��E?�{�\�q�R�����`<Ȟ����R#7���:E��
>�1�Z�-�4g���c���7�~al!>a�g"��f����r2޾��C0]xH�5�A��2^��n���E�3�.����n���������w�pKw���E��f�т��wA��P�F�B�M�x&����fw�{Fި��Ә�.����M&$B�D��[��������;�;���u���Q��݌���Tذa�|�p���;���=�h��15�ɄL@� cA�֙��,�GiD��u.� �C�b���%u�(��C�ژL&n`mk�R�%2#�u��g��/D�x"q�^��i���w�x{pJ���+}���������ݠ�ر�Zc�HT#�qՎ�O�cF��w�íN�<N�8։t�ZJz3j�od^��~�v.�|b�zk8ʊ�*Àb&�u[fJ��l��ϓׄ��x>癸�1��nO�Ȋ^V6�yG�7ފ�f��]�L�x�v*��}k�H���yPژ�v�~�F����(#8״����>oM���n���4'�t2p��䕃����ެ����FH���t7dS#�{��1�1n�\9�WS5Y�XE�p������ �3 у��c�F�T�g5,b�&O��b��FD%�s��<�6�Ρ�:�lY�.f�(�z8y���)'�Wⳃ��b�I��lZ�e�9xPj�׷��X�0f��@0�pT8C���PQP
��׃��������ʹ�b��$xz�2�rx���S�R$`Q�D�4��i�U��%�Q����	s��[��p�}&�B����\tO������M�Qs�`�wу�:����Vi�s]X6.�]�G��x�e��8I��b�kФ7���F��w{��~�(fO���}��Z�[`�y�3�F��¡�;���D��7�7-Z���:�t=���xP�e�0(]*V����i�6�ƛ��m��h�8�$B
˰�	�D�������GyxW'BHm$$XЉ ;�?5g��n��c By�� 'Hd�"�Dd��1B~VI$��vQ0C�Bv���x��HrҤI��H�Y$�m I1��oM!!�$����	��Bi		&$�$�O�i&�>�c0�ĭ%X�W+H�W�5>B1� �,�l��4~��u�����XmbҲ �����d<�߬�~�_��}Z�²{}�?E�K�~�u~ݽ�$��e0�zx�<���0�,��j���u��b̢k����z/;�&%�*�I!�
�[�It#�k�-L�I�-D�H@����� H@���Ap���.2<Λ�V��TPjH�l�/�D���d��9�~�VCn<�I������O�$�δ�ӽ�P�ԋ�ɉt���l�$��(:F6Z����RZ���AY\�r�Xg����A�}�/���c\IH������ HAd�@�!1?a!��$"	 A$ �H$�!�� I �d Ȅ�I��� H),$�Ւ HJP��H� ��# ��	���$	!�@��A�&~�f���K�X�P��)��l��y���^bA T�(W*�5�Mg���%w�lH��Hy�s14�V���F){�)ގQ��̔W�v��y�H�QQB3ÐjP�z8W�>Żp��������7f*�H;��v�k_�T:��`�[�׾d�,���;��,.�s�$��f������q��Q�Ȇ3�RR�힂��ˋ�L8T4B4�  �I�h I!�λ�4�6?�b�0�pJIH&+�!*�H "b]��$�B��~����I�߸jp�=T  �8�9)��p����Lx_32R��W�K%�� �CF�Nrk&�!������O��?��I�����r�ꩭ HA���ؒfŤ�D�	�0�Q��|�/�����y-a0�Q�W��b֘���={cj�I%��]M$�ɸ�&�* HA���Ka��.�α,�r
�4���(���`��7���0p92iy�߼�v��%jia�t�>[w
y����	�D�<�,
�T0ūv� �B
���i2$�*���L�t\�)��j�=sఒ�Y�n��L�W�y�B�R�`O��,�@$ ���q�C�^@�l*�,�� m�"F�rk�T�W3���j��r�X1��d�:�@���P�N��ѬYb�H�
�_{�