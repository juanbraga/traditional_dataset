BZh91AY&SY���� .߀Px�׿�߰����P���[Se$�)�����SO)��A<��F��� ������#M���A�LMH�!F��fSje='���1Ohɉ�	���0 �`�0�%4��y'ꞓ�   � 	G�
�"D�\!>�滼>�%���2�?4p���,����4k��kݣ,��E˨�u�o��S��e�g4�o�7�ӄ)*N#ù��$ms�}57���o�;JHU��d�؇%�4�}3�������}�5�ծ�k�30�u�#)$��)�:����6�Kl`c�^�UI*�ɑH�~H�bM����}�~Γkllm�m�A�_�OL���b���)6e=�ͭ߄��c<hAL>��Bޘ�G3*C�Q�
�f�г��vx3}��Q��� �s�'�I�U�����*�5& ����14׏��*t�pøw��]���JS�j���c �,-�ʩ��G�Q���~��r���F�հ�X�$�T�0L��"�#����8�K���
���������
�Ubp��e��n�XQ���W�c�a�j�t+NS���}�eF�H�x��T�L��j2G���(��q��U)�{�c-�6�p�	Q
��-��zH��t/���A9g�g�Q�=�E���n�r?T�q���T\B���T�33Ԡyf��9�jV�����2�Y���9��	�.
L�
�yq�v
�%�A�ə<2�v^B����SHQ=:
X��]�ʁ)2�;��&0��2̩w/ ɢa�g�H�"�PW����	n�!]YJ��t@=����w�£�Ƽ,݈���r��6V0��l%�K4����5�V��E��=�U#Z�՝��8qJk��G��gVt\b~9�X�	�;���xD���k���' U[<��Hצ��[
����e �2�w$I����,8�-E*�����0��2T*�E�����ٗ��B{���N�A�ɐeu|m��.�p�!�[q�