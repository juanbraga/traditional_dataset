BZh91AY&SY���< 3߀Px����߰����`�z�����{�X��I���S�dɢ�����4 h��H�U !���`aM0�L�6A@�����14Ѡ4��S�`����4� �c�0L@0	�h�h`ba"!4��M�I�P)���SG��#&��19RU��HHPE�������+,����#����#��f �Gk(�b,��tp\���n��F�!�"��6�o\�B��J3��6^Π�GD�pW
|iR�%�&8$Q�1B�Z�M��//E�uiL�&�;�Y�z�BFo�y�����$fp3]�0�O]+�A�*�% ��l��-B��-����/��͡�/�R��r6<�G��Aő��ɠ��̋�%��B�T�u��͈��Ѱij�v]�YmjY��� N%��F�L�l��J�}9lm�"�bRr����2ڼV�!��`Ne�BP�X�l�Bm�U%s7/s�YaR�A�BJ@w�_���^f_�}a$�3C�Ν�����W���g~[���ea�Z-��k(�@�;sn�e��
D-�t�����"X6n�@9�l����H�d��VA��v#m=�v�K̭`3y���x�j|�gA�U��%�ˬ�	t혜��G��5ltx�vX��À����3�t�U�`�Y:���>1��A ��$��$�����S�K���u�T���H�%�r^�G�[H��P���Bɵ�#esQ���+ �� �Ide�ݴ�(�(�g��p �����5��ky������W�%՝/��IX��.+@^��c�9e"�"�/*x=ȁm$h�����c��c�@�1�����ȼ���c2H��1�
`虻3�{I]��*���È�/�rݚ(���:��E�B6�c^�����3/�ь]�ފ�1�8P��bF��H���MV�F�S,Zԑ}�:���척u��n�օDV��m/J�FE|�U��a�벡�����1 �%��0��5�:�	1���`u��&E ���$����5x[����<=;�r�_lp�d�%�A2݀��K�vZ���H	)�lPQ��^��["�h�N�V�N���J 5�ά�H�m�7c�T��ڥ��
�E�3&8��1��O��O|�ݬ��+8�I��ʄ��]�g���W�P1O�苏�a҂���c y��J��!�8U��a(:���mJp��(�Q%����U�2he�GqĲHEA¼�ov	ɶ��oB����6�3�WY�=���冰��[셉�r���Y��Z�E���9���}Ѐ~L� �L��7��@���5QS��-˫�<��f�!�r՚���9�[�U�h;1/}TmS���jGf�"r�QiR�,��಩�M_T .1�do��֋���0j&Z.4�:�멥���j�D(��n�X/�Ҳ�_R��kJ{�kUJ�#ef:�ѩ�R�)���;m�cl #�&�yi�X�ܑN$?e{ 