BZh91AY&SY���' �_�Px����߰����P�sl��:�i���F�beM�yM)�����4��� %@       JdB�D��M#M=@  �	���dɓ#	�i�F& ��j�MO4G�hd�4 &M0� k�J-�����������N�a�?t�tPp [ ����D]��:�]h�2.����y��v�Iƥ]���\��Fl�pȲ��k���T�V�����q	9P�rg)%q �8��W���!j�AT�sLD2�=��N���t(�1���v�_u�pq�'1����ޛo�M��ո��сo
���,�b�1�y����ԙ*.�h��
�6����4.
S�HuKs������&�D�gA U��g)�i(L��f���d@����`!�A�I&!�%���� �%�e��I�V�F���IFIn�b�	�0��"9H	�ɚ��&d�r@v ;T�FX���8�BBKbHD	��έ$���Er�u:���5ɛ�a��MS�C��E�	��x��M[&d�(�O�Up�$U��w�ph�E4�/ɼ�?·f��������I1�,}|�2^D���r�,�Cգ0�B4q��]�zKI�Cȁ#�wT��}��A����u�=�Ô�N�y(��Jm�$��W��`\�$#�s��]��LF��>OE�X	H܂���g>|D����̳���3F���&/sv�����PD=CC��g�(:&H'L���V��D�tn��^B]gN�L�q3_͜�0|�&<�4h��p&�V��lxY4�e��un�*d%幐2�Ѿd2�B��<ĥ�'5/���\$"�1c3&�4�v�RR�k��q�NS�rcZ�˴�2���h�Q�uNA��uf
$�ĝJ�a���k*!���eBp�[���B�aMʘD�0��Qs�X��@�`����c�#-��!dA��YRP�Ϥ��s�$�,�	iq~�F`Ҭd��:��R�!m��� �H�a����Q$��T���8oi��8�)P��d65�=�Po��
�đ���IAJ��7�R+��~����ꨖ1��411Ka�aR�n�ͫU��By�`^��TZ�Bƣ�0c&r+��"r��p�(fZ����-�c�}&�Kq�ɒ�j�����ܑN$'��I�