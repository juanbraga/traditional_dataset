BZh91AY&SYg��[ ߀Px����߰����P�v�qfcHP�A44L���=	�i4�z@��A��2    h   $BI= &�=�i�A�Ɇ�F�h�M0���a2dɑ��4�# C �B��S��l��M�S�yM�h�)$�{{�v$R��HP$���������oHCP�y���i��9�Cv�k��_�F�7q��ۆ�"ܛHo���pq�8Pϡ={ʻOQ��Tr������Q5�I�C��{Ԏ�Nk�ٓ����	�e3e��op��	��6���Qnt��H���A �����$'`q���|�4�!�4��#m��ަ�_w��L/T$-1���M�6A��A��NO���k�J�� ҪkM��b��՝10a��v��2Β�C����)C *�N�E'���V$��kG$�*	/��D�a��b����tE��R�`-�Hx�J�
�vI�P�v��@i�K�.��Tֶ:��4�\͖t,i:$ͩZ��T��N�E�)�����Z(�٦*p�F�,���2�ty�F����1���DOV�%;�h��Rʱf]W~�8e3��gY4�G�&q-��gᙰ��P�ڸ�=�$L�{����-��6��\=���&ō{)��W_cjl����x�+]�{������==�:O�����g-z������{��<�4O_��Ā�ɓzʾ��}7��� �(BG�l��A�C�b��EyQ@L��B?D n��V_=�FdI,�Q�^��Ȅ�.�v��P.du$"��G&p��-j����WNz�F�`������sߢ�'3����s�TӨ�n~v���,8��Ts>���!�!����I:P����T�}	0���!����ځ �R��&RN����y ���e�г��]\Y@L�U��D ?��lt�5�&SȄ�	+�գt�R�[����4z�O�
�7�S��b���&��mA�(�],o�c�!��2a������7
?��	����W8.5=�l��x����;O�������:F���HΕ������+6����[׮�PsJ��N��Dn��E��Ë+�d�@M�"�.�t�"�&�xԐ�sB.HF��7��"^�yci>j�����I�hOA2�9�-����s��26�J���!�^���pF���Z	���SQ;I�YQv2�fJa�%�E� ����� �Xz���)e<e1��)�RXE���c ��T�	����6--E�8!X��J�Fj�]���z��}d����\gK�Z��޸�,��=MZ�c���.�X�8�T�2���_&��D�6��{�;B�w$S�	{%�