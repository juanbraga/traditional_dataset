BZh91AY&SYRX� +߀Px����߰����`_/p wI
T	$L�lF�LI�h���L�24�4"x�R��� ��C@ ���&L�20�&�db``��4DF��h@    0&&�	�&L�&	���Q�L�M�)�J��6���z�P�=L�T��#h�"��.�"ǁ��J���R�!�0L>'�X��U*F ������AT7�OE�V��鯦/tܭ�^q�YU�L�Bë�[5�;+]�+;kB@�&�a�hPJ�m! sr��P��*�@%Z?̻�(wӺI�X���W.5B!�4�1��:��f/��(Z��"I݈l�7��o�H̙3[,6)����[��gu�Iw�G����w����)9ِ���)1o���y�[c¢i�7����Ӯ�\��2�^4F�Q���t[�3t97\R×=�� ����'lꋹ"��t���mV������F賳�+LƔ)�r5�P�F#���(Κ��؆�2��dr�����(k�o�z���4)��W���nӼc��b�kt� �e�KГGu�J!�C��Bz��.�뗫"��X0�9��;F��5�=Zh�M��,F�D�7uE���*8� L�S��uR7�:�"]�\Υ�p�����:O�{24Q�0[͆��mm�$*݈*��{|눝��V"�s�����Z` @p�		I)AO���tP}�U.X��Z^
Ǯ�)p<`-�0��Q��I����$�D��3u���Ų�`-xm�x�J��!7+ t����l8=�t�]���Ǟ����J};q�F
) ��+���NKA���n�/	�L4��X|����7 ����(�y۷S�r{��B����{��d�?)˱*��y�U�搰�J��|�1ǹ@����vn*-b�b�&�{��	̳Eulj��lka�%�h�#��F��L�/�=��c�9oS������Y M8�-q���O��'Q�r���1:�p��������Q�|~��gA�(�s�|����C�8Q@os�F
9��-qΧϋ]���'#ʢ"7]y�d.0fā�b��8jk��C!x�
FVfL5�3�O�����n4:d4��EF7(i�z�`���`z=4�����pǅ$lT4U��*�F���,YTd3`���«%��(İw�=6C ���"l^��!K�!��XJ�`g��x���\�ڠ;��\zvfů�jʶD<��Po�FT�LJ��z���edq�K�@�X!@co7H�)�zM���TZZlcsI�.��*���8��7��V�J�jά���-
���z����0Nd%3B���l�(���2�6����Rj�C(4�:�(����5L?-��#�d�
���y�oX�qV�W*�m{�i��_��df\�
�]I��md�5U�m?�w$S�	%�� 