BZh91AY&SYۚ�� �߀Px����߰����Ps���B䐱� �@�M4ɠޔy��Hш1����h      BD�OBd�4�A�   �`LM&L�LM2100���zF��Q�i�ښh2�h1=M���]��W$�JA� �gQ��y��CTب���v��(�ɍ���2����c|���ϭ~"HC����B��4��H���蓋#��g�@�|}_���!L�!��I �@�6�r�U�m�r�.ִNW���&�f�b�\ٱ�s8���k!�i���;�f���H�l��/���i���X&�j��ɰ���"�#خ���~M�co�/���͎,���z�l~�>b�&&�R@D�� ���לR��&�k�lI{e˨��<�a�Z�K
�o@ A3�v$�u�-��ҕ��J2�f
��3�C�
��x.4��Po��k���7g��1�Cݯq��l��ۨ�/SЧ�ʋKF�QZ��|���oG~�#-�AnDof�2�)J��D��2���#;q���%wdU%��E�h��b���̽%*��J�>g9��ֻ�S���i�jB�Hj)#B��-�܉8��ϛ��;M�����l	82�>�^t������`�J�%�O��� ���.f�mT�I�ht��˿sQ���$���a��<6��l�-_�����o6j���w��t'�4�����98/�ϓ#G�1�}`��#?���D�����M�}Vp�Q�n���z�����}dvm�9�xؕ<�Og�i������/�y�fW�aݖm����L��$��]H����ٮo�8gK.�S~�[簆�����*9|C��^�,�2�t��#�.�/����c���ɮ{�*�ꢡd����ķ��O��0�4_ɳ7�@f*"a�:R����bŖ��Qo-8�b�5���V8�@$�3�Fv9Ll'E���w�0�d-�x1����A�lҏ���������S� ��r���,�ٴqxݳ'�d_Q8�fJK� ��"i,u�T֭��Ҵ�$*��fL5�n��:o)�?���ceG,�xo*>�'�w)0�G^�]A`���M-�#++;o��4P���Ehh ��q�W��|�9�oQ"�r&{b"���]aˬ�V���{�<FH��3A�w�@��t���$.�Ir�q�&�aW	߽}��:Np���Ҩ��m7x���^�0��Fx9m����Q�B�I�h|a�	J�:�1#��M��Ia�5��q���I�Qk��1C�|�a���h�NʬI�=�k�(,"��jKl2�O�Um��R��@��2pB��*l�d�����]md�]&H�"x�[fA#�f�d[�vS��l�_W��F����hX̏����UG�? �u9��3&A��W[��]��BCnjN�