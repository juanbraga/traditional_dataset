BZh91AY&SY��z@ �߀Px����߰����Pxi!����ܵrxI$j���J���꟩�<�S��yG��i聧��I@�*=jz�P�z@��   H�A�a�CP�C@h�OH`�1 �&	�!��L����S��24m �Phhh   �s�*Љ P��B!	�K�ߍIbF�&\ֳ���!�J�m�����{����f��Ǧ�<&$�9�DY��o;�7�f]S��5����2��Y*F����a�<`l�F3ޖiV@Nz��ụ�m�k���&ƛ�n�,i_�����w��#��[��{��,5]�*sN�~��-b�b�s�,<��M�C�V:�3M�7�$D!�\�g(^��Ni�N3D�i��)2��+0�U��!�\��t�L-���W5eB����z9�6����m�p2{n�N�G/�����Rl�=V&l��{��N�BX����8ꘘ2DJw2��u�0eZ�U�6x`Cb������펗wA}��˻f�c�]�9���_����먑�2�:���G��;xƸS`��7ǧO�Ә�h��1���;j/ �/2�J��:O�8ԨCh^�/���Rbu�/�D��3��pN.�x��h�ԅ�1#�+b������L�����ޔ��"�*�9e�ݓoV�i�0�"�����p�n��!B�P�L!B,3�O�cc�uPZ%�B�3dI�����������y��u�냇ۃ�	��Q	�d���]��OV�-U����@���fp'���
�jp�*_o�RX �c3&���+�d�c���9L%q $_0!ql����',�,�b�U�CīQS0Q<�ԑ!��/��aJL��H��ΨP��,��K�T��#%3B-Lc- ��O��ި�˦�J�GI ǘ��
od����m��ܣ�pKs���Fa���L�X\ԥ�ܙ�PҪH6E��.7!9l{�\�Me�"dj�*P�E}|�އ��ϴ�-W�ll*`��B���4��Ѫ�E)�ͦ���f�Oš�4d��Yi�Į�*'&�D�d�#'�9���,*)�o0�NDs*U�Ee���x�f_#�>WH��kd�cGvH�'!w$S�	�7� 