BZh91AY&SY��" c_�Py����߰����`x�n���>u��ju�i��� �i��5=&��x��z!�� MHh4d�h  Ѡ��OҐh       $Ԓb�56D��= hi�P�F��!Q��&4�20Fjhh�FA���
i����S5?DA��� �h&��}�#hA�
����4��:x�fI�L1P'D�S?K��縒M��/bɕ.K!/Ck��[n]�{�Y�#jTX��P�US\XA�Ds��Ǔ����՛A��wo�ᅝ¬9�r+CT�6�\Qxg��ǁ�������D�ϝ�J��
#��>l�4z,n�/$�f�|_A 1b��S+���)2��	5�������b�3!�+��(|��3>��D�!v2+q��c:6k%��R�M��L�H���N�������)J�"�2�(���fC�u\KVS�����;�NF��] <�I��5ɽԴU�^�f��1��+spF���G|��FF'G������j6��jٿf����ƭ�_-k�:媎�)"F���i������K�e�Y#�2��`T��y�`\�,�Jm5A����T(����"�Au0E/9�%l*%&G�t�G/dy�E�b�hK����me��{�R(N��$���PV(Se	�4؄Uf*
�6�rdI[()ER�xF fBlBnW���5VL(1e����a���*���~Ɨ�M%t��ߌ�qt�ѮP��	:Y�h�o|�ާ=������������T_�����~9�㫏��kle�<��}���ϊ!Yk�X4Q��_A�9a��n�!�D��E���7�S�y�6��)L�
a�L����R\�n��*s�i�IQ�L���J��u��ӹ�!FR0d�_�H�=��y���i��Ӫ�҃2��%G^���bJx��L��I�l����G�^�N��{��U S����8Udŭ"�/��k�6�ƛK̅���A"w6љ��1*9\M=����*�PKA�$�l6���'$A�[��K��`j`L ��ɥ酵'e�9�	ݬ����@X�GB�8Ȍ(�(�.�k�!��"�g៖KL�$Tfa�2l��4��L����2�c>t��V��AJ�J���+@�lAs��%Z�w"
i�%?0J�߾EZ���%��hR�Uf���s����ya�Yb�����N,�6�Ɣ*�٤�"t	���pi��,��*�ܷ�[؋&��������
��2*�C!O�Dym� o����Q*K���0s+�I��sj\D��R5_��Ԃq$6�S�4IT�:��Ǜ�b��y���oL�n&4�^�n���{QvAE�й�{5m�6�_1�(�����B�ÕDT�?��@�ˢH�����;�����2p���d��)�jVrd������hI5�9���Mx0)�C	pSʕ��z�7���M+��̥��ϥ�f9�r�z���B����)����