BZh91AY&SYbb(� �߀Px����߰����P|�{��G��5�;:�IdɄ�e2zF�'�� h5O��=@�  4    "	I�L	���`0���C�"M����i�	��d=OS�zA$M!��O�x�S4��1&�F�� P@#p*�I� ��?�{���p!�U�P�2�$�X4���7YG,3����ݗ��KVS�!���a��M4�"�3k�+kbԊl�T�*:���g�4:*�;�2-87~B��!02�w�R�HfUotd�0!��	Y<�����/c���
�CF��m��V����]-X�����3�:�X���"7ɺ���u Ø8N�6��͠:jh�3l���4Ă��I�-h�I�ٶ�aU�!��.cF�I&��d���v��{�у��SU�cuE�COEĠ*��[@��-��ӆ�8�f��3."�6D!�zZ�����nͫ�����p�yo���T5�`�T�f��-�룻s�4K:�����F�$�IJ��Bů�s��m����6 �ޮ������B�Hֵ&̣ٱ3`<�Xa
����Х����aG1�t�L=�8u�FSUj̟�Y��`czX����wcCq�����+�˻��/���Q9�a��7�
	$�՗��z� �gl����5�����-��(H& �`��Ջ��}����ѳ��H�W)(����u�����p%�L,���1L8�����*�GA ��Ȥ��Q����ܺ��̴�q���I'T�0�(zu1�rC�:�9.Sm��s8-�	�GobQ!O0�y�:�H�0H"��*ZC%�I$΂��&���i���˕�aF눃�B�aNW& �V��t�Z�.&�DQ��|q�Jf�yPV��Q��LeW�<���8j+~>�$��̘k"�p�ۇ�wL�~F������6t�^���`�j,5�(
&ʴ�`�i8�@R���C���U�Ɉ@�3��%�q������gLv�}3����f��%2h�&�-X�* "��k��b���cM�$�I%�L-v��J�_YO��4��1�8S��ٌ��Z�1�����2I&��0N$�>F d��&��ͬ�x��mn�l�OJ{�C��ˉ^�%R�f��$�}J-NF$j �!\`Vw�o�6��e24$���I5Y������pP�Dp�V�q��JIn�	���(چZ�ɡn\tl'ҩZ\��W8�� �K�9��=?*6�Y0+����)�GP