BZh91AY&SY�� U_�Px����߰����P[Ѯ�Fm�feHI!4����z��#�dѡ��Ѡ�� ��A� d   ��"iG��)��h z�SOI��	���dɓ#	�i�F& �"Bj� ��S�#��h 2 z!)	d΄�Z(��Oi�u����BLH�L�\����������rҳ/z����e�Z$��-�sӅ�c��5�2����	q�8�C��J2����CS1^�����(o���
� ��2���mJD��B�A�$H7�p��f�2`li��]����c��� �F:�q�rSLR4�б�/f���H,+p�ϋ�P�B��at�74��K@�2`B��00�!	i��VdJY;������7�
%1�C1�G:�B�e٩C3$zigR�5!��B�!���5/h�Y�b#(&����V��[�L;#:*��!+�d�D���vR�b�b������o(v*�I�H��H�#q�APY��uOm{�i�on��im���;l����y�_BlV'��2��bf�-�/e�p�B�b���h2�X��arp�0eZ�U�[�p��mlW3�u;��n#<��_�m�׿']�������x^VPwUN�g&�T� ����}��z��ݚ�~�P<l��ik��q�m$n�ȁ/!�U�Y׺-����P��%��d97���[i��j �����b�N��`�@]~S�Z��߉q���,\��Lq���ӱ�^����P�3��￘���Zy&g��=ԁ�M �H��ȅ;d\�o�+�a�.2b�	8�b&�nQ�v�?W�kd��S������gʻ\SF��@%J(T3Z�*ql�l��F2fhN�e�Q81�*1�b�Lf,w
pҲn��� ��m1��Y٠��*1�|+Ͳ� b\��2BZ�o�&�Q`Cĕ�S�Dx����\����k(�a$A	�f�Q�R��nqR��(	��W#���'" �K��s��p�c�	e-d����
�i�=7FA���
w<�w���I�F�φf*͛ �N3p�86�.�k���H(A麤����Q���QF5��s�,� g�=�:�>�r�j�(�� 悉a&Pt��q����T/��S`$�OJzfe2�+P3!B���E�a*����l��P�N�ǡj,Y���3^r<�ILʵk�i��ƌ���v)��c�Q�I����=��w$S�	��P