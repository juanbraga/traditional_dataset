BZh91AY&SY�$�� �߀py���������`_|}�=�{����x���hTD���F�zh�j=OP���C� �4h� �2h�@h 4   ��db0�`!�M0�!�F��i� �ɩ��i�F�OS�#M h@E2�OS�ɐhmCM� �@ 4hHD�2i�F��������ڇ��M2�T`�hU��$� �_��$��T����u?�p�"ʢ1��e�yA�uU�A!">^�Cb<{O�{�D��J�H@n@�%"I�B B� 첗�I@���D�$%�[��<'�����0"�Fɉ�Z�H��cl�J���.�	�dIa-$$&Y�avtSN�BrS���w^=�<oDGt$�ZNs���g�gY�� 0�s�,'�&¢�TB�4"j3�GsYTM�ů�ţhZ�ЉT×6�Js�Vܡ����?�����s���n٩�;�b�~���&�#L��o5N��xK�*C��r8)<<-���%3zC�2�32�)s�&����#p��-�|9X���n3rk����Z�d4C��f��I�bL[5��8[
�zL<i���Ӽ�!�a+z#Z�.ctbv3��P�:O0`���KS�>���y�3�k��Lq)�ai�XJ��8xq�Kne��)�� ��3��sCM�C+2hĹ������ٝ�TvN٩����P���.�<�my��h�,�s���)�m�S:�*��:�Vf�%�\�Q^ֽ�k �1ܥ4b��N�ŕ�jWӅ떭Y�J%t�-1�1���t��U �T�M�㮴]-�C�F4�]�I�5Rz���Ma;hpV��f3rk/�̌;�8	&�/V��iD�[.7BSDB���_���vmt;=nӉ���QM��ѽ�t���6Ծ:5B���5Q��y���:��۳���| YݒM�H�D/������Q�iR&܎vBnG��e� ���2G*��Dr���)/�[$V����I*��q1L�@/ayb�'���2T��������	X��%���jyJ�g��dX] 9�<. ���d->꾔$K/��ѻ���#�>���X��+ґ������ǖ�a)|�p��>�ԡ��}{��xk�3bA( ���Cvd�p{�^��Muݢ�]	�>#(HVO��sqe]�TԚ�R�Ե��P\wʿI7^Q�������Qu�1>�~�F�脋�0��@�4��M��FP
19)���=|#L�궄�1�,�ݚw=��:ͥ0߽���2l�b�I,�=	r��YB�9
��\�X�p���/+ޖ(�v2�"<L�%���������p�ĳ7�X��T��	vL{�o
��J'pum���[�~��p�(֧`D�I(�d���.M�| ��p:�J\�%;�f��<�k+15P��8�E��5�BJt�7��r��/��><�{,J~��,�x6��3P:�PuD|i��nLT���h���U��rA�Ax��%�F�	��L�V'��H�2G�� w��Fdl��Jӑ��T���%�R�))0d�)����Yd�����ɀ�m�c��QGid7%M U�^C'e�����Az�Q���H�a4;��7q��X�T���v��} ���:�x)�B��Sc�r�IDd��n>�𿣓 ���3�bq�L��ARI.�:�U'@)�ݸ�4Иt�|96��J��7T09
�"�K;�.1+��HB�`�H��a�f&Md�D���ϟ�\���d�4�F%I�������؊�=# Yqٴ͊RX�д���綋Y�y���,U��}C]�Y2\����w$S�	K* 