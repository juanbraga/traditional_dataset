BZh91AY&SY�b �_�py���������`^=/;��|+�}Oj�l�-m�BI�@$��M&�F�2hd=M ��T��))�       �O�Х�5�  �M   ��"	F� SG��h�  �$�T�SiF&��4 � dhh"�Bh��O�1SmS�'���SOH  h�F� ��[�P �x��I% ��'!������0$ 9TF4��8��NK��<�8�D|P	+�;����v�4j萵Y	� HU4��hB�!I�w1RR����h��&��{%�i>�lLq^	ĵ%l�Z�U�P��C�l�VeZ��<3Ji�I�	�&K�L��'fN`������"�I��+'V�ELFwk9US�<b�^Wh��F�)-i�Ǚ�sT�G�eQ4���ţh\hD�4�Ѯb����A����?l0��e;�v�ʇ��pIڐHIb��FZ��t���Pӄ^��UyR��cD%��T�e��}d����v;��ɹ�F��DF(r�<���^Sm����'a��94��EGFh\&	���}
YW�<!�Vg:(zf
�J�j�wP��Ր��\��p�v �F�ؤ��`��Ɖ���Ar��*�B�B�5���-��OJS�A�z3sF�&䡖�7w'h�\�EF�B`,c�+�Z�p
*�)������,]Y���D�m�')-�ʳ%N��L�[f����
��Q���m���7�w�V��G�T���C�Di��"��ʅ	1k���.�*W �:6��T����ֵ���*�V@��W4"{ˉ��LDR쁝��L��-����%]�r�*d0�
�$:��xW�Iz�{58wD�^R��eI+�R�0�ndP�1&e�3d�uK��,b�x��ߓn�Io�� @t�
4Q6���F(�f]�<�m��y&ӈ�Qk��] ����o1�
-PD�9��+>��E�����`�4E ��勀:��e��X�G8��0�8�l�c_��Tˠ�UU���\�:R8� ����}?H$ݗt�����İ�vW����G*ґ�oO��u���|�Gd{����Ā����1��6�b�P���k�$���|�ڀ�^���.fQ$Q��H�<�A��6��M��,�+�JT��
����M��0tl�9�u����C���M��#���:��At�}zs�T�J���`����O+�$���х�R��&�>�.�Z�i�j�{��$�D���*�j*k��
֑"��Z�P�Y0-�K�����:>�Ĩ� ��fd��a�e�+��Ed"Oً�1XD����HEvTA��xKo��5d�g*��r(M�J��k�җ�R��u�u��A	_Nf��A����&ca�Wf���kdz�W�F�Ґ�^�Ɇ~���o��i��rxA���������oQ�=��)���;x�5H�������PlT^`c�sq�n a$�%;7�-X���N:�2���6̠!來8 jj\�Œة{�^��[������Q��F$�♄#~��qآ>���fb&	El��|4/wt��E&~gn$=�ғ1կˁ��@�!�r;���°B�͍M:Uvԅ��n�.٬�F��F]���S�ub4k��0H*8��eʆ��j͑[%*c����tMI��Ss�7ᠨM����e�`���\���$�h$!Pf�,�lh//E�8!c��+���mVC�<* M�k dgԟC/IT��>2wx��]�t9��-���ꅬ�9L������#.r�� qНڀ��rE8P��b