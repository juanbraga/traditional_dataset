BZh91AY&SY1��2 1_�px����߰���� P�weg�����Q"OjzCSOF��$i����FF���J�dj�H�       �Є��������RzCOPѠ  4h2dɈ��	�����$H�$4)���2z# =F#I��
Z!$��'��_�ɝ�T�h�k��M�~�
рR����4�[��qy8/�[t�����yK,�xU�ޡ�;pt绠M�lz�@tşҲJL8Y��[�N���@�������-GMa�V��������R�[�5��f}�K2�\�e�2C[�Yv�=/��m+�]uBGG,���'���T�>c���Ym�u�\\Tu����jm���Sm�j0�6�*&�䒥
G�U�բ+_��x�����xn�V�M@N�{�ADMN�ڒ�T\���d���x_̗Xv`���t����Z��^�2�Eފ9�i7�"�w�:�Ԭ��~��!�l�kŧ>j��%B@ؒ�Vd�՜�~�G�)B���b���ېF�K�d׋1 �&TV�`>&��&�IDMى��S��Xbe"�I (�s>z,N�R����\��
�3�u�Ű���ɋW��;�w��rZ��C�:�;$Z�[4�\�KϽ8��*���E�	TB-ϩ�X�s,PEZ✧_h"q�C d��\IfNt��w�L��R��n9��k��g4���9�`�3�_�8~�۪k/Ғd.�6���#d��)R��D�B�l9b���95'�E��p>�0!��@]-8������H�
��p�	$���!8L�B���+��Ь"Yȫ�j���Ag����[;X�.�$��{���H8b����#v&e�0��@ɘ���L�A9&%�2N�h�!5!�q���9��z�V#a~�T�z2���1;�J��Q���xVP���f�B��,�`<&�r5�(�`���$�d�.�S�Kz�LV��&xŉg�$_��F-e��,J6!,lKr�UM�Jq���xxD���H�
6��@