BZh91AY&SY���^ :_�Px����߰����  Pl���Wn�a�SѦI���6�1Q�щ�C@��4	BLL�S@4��M     "SS�hz��cF�A�� 4 ���L�1�2`� 4a���b��4���!�  �̀�$A ��@��9Ggʧ[J怨�k�检�,Ff6�3(堳2%t�쏗/����R��!��> ��aX�f�qZ�׫dp��*�)0�f�3&Bp(��U�QV��H1G� �n���񍦛՞��Y�U<��Q�\��F��5�5��P��6�������S
aܪ+Q6q�z�Vօ`f��jB���xu�������lp3*y6���RѦ����jM�G�e3k1|�.��g�{C�؋J:�T����Fj�3;ɢ:aAf%e�VTg8�7;�v�W�֣��h��}cЌ�8p�&�_��r],,�^��:�$*�Ϣ��(]mQY@�5��{�x)z{�?dvw��Cc���ߜ�mT+�Bɱ���u� �~��@���u���>p�13��eb@�x8�18kf�ץ�ޅ$�i�]��WMh�T��|����J���HzD�S	1a�kK��o��Z��vAA>S�)�e򆵨���}e2����n�u����F'Ȇ��G���f�����)͏i�#$�hL�s�@n˧��ZfVkm�<���:�UH�sZ���h����#Y�y����|(Fb�st#"�g<��QcEM�$@w���dĠ&�����)�E8&r@F�P^�u����ɢ�mՎ2�
��|T�3T�!���J�Dڢn6p�*�Y�]�m`�3��.�*"�<s�%�2*ɀ�e��g�������ӊQ*QRh�5���N������8�^�N��x�*�AIi\�쁣UȄ�[�"*�F�B�QQ�jZA):��ʪ�/��&�Aq�V��%�b��; mSB��SiG=3"Qp��
*B ^�k��H�rE8P����^