BZh91AY&SYa��- X_�Px����߰����P8y3��r	I�Ѣiꌙ��7�M240�=C@�L���&��4�h  i��  DBLD5=&�f�G��@�M`LM&L�LM2100	" �4ɢ��~I���j2 ���04�$E�P$������ҳ@u�!�����A,f6������dz�m�f�]W��",����}䶼"�_#8�6���G�na
J��xv8W��1^B��i�*-,�JY+�H(G]~ͳ����!����2fxܨ��x7+w��|���.�YD�ţUP�4���Ɯ�J��b��&�/ $��2�(Xp��.d�$���C�8�LU�W����8[cco���48:��S�(��B�Ug��2���f�O��)e��T����1	v���t�/aV�^Si�m�i�2��M+��s��y�ݵ�0�V~�ڶI�[����h�Jrγ1���?k|)�u��*0]x�M��-�i�+������yxJ��'�Nw2i�E�#�06�1�*}g�s��s�")VqON���FcV�1�^%��#�����%�L(8�t�q�L�N���n��3��_E8�\Ӈ�&�wNui�p��ٞ9�M�����!B��a� ٨��T\q��������U��S)�%��]ϻ�=�!l)y���NG����9&�d�80F)�
H�I63Z��Z�g�d�0sRJ#�m�&�1����b�ԜfjB����p1�����%�H����J�C@�M�3��7��Y�,�����!�6@ҭc��$.���Q<�Ԑ2vb�JL��D�&tB���2��K�T��&�	�KVY���2���.�2�'��F�V��H�F�����;2͡8��r���X��n4_��4X����-��3������$rA�s���-υ�(#lʝ��Y���f�2!�E;Tv�]3`�jn#3�xKQ�Pe{�ef��D+J�Nŀ<e�ʪ�Q
*8K
ѩ9H-��M7�^�a�v%A!�4�����U����I�V򘪕n���:�}L��\��s�|# vL�*}���rE8P�a��-