BZh91AY&SYp�~# @_�Px����߰����P^�]�
�Y��H�z4#T�?��OiC�Sj=G���z��4�M=4L��412hd 0L�DAi4��DhzM=M   d�s F	�0M`�L$����4i6���T�Rz�S�4z�0@ =M,��*ĉ@"�I��r��P��Y�:FC]"�Q��!�Y��S(堫X>�Q��,z:q�Q!�wr��$��@i�Ba�?Y��3G`�h�%Lv�K��PH��%I�f�5���!)d��eG=a��zL9���&hwU�p���=�s��IZ^vW蜸lq;�1�nOO���F1U���/WU����UT&�su
��ryή-f�����m�8=7�S�E��}��Y/�#���d��KP�ŉi�b[$�ы��C�Q�
��O��ĆX��ow.��:�QU[ew#�ƃ}�k������pG)���B 0��igB�R��$��(o�c:to�8�R�=��e4���e���������J!����ÜS3Z�6�؊���B*V�\�.ֻ�/���O`X�b⅌HZ�ڽ3
�M�n�ѡ�}�aE&W�c�Ì���+FSG��]��2���	;P������2F�2�� ��T��ԖC�zw#@ǲb_m
���p��
��ڀe(�i�+�M�m�V��-U$��dPG�B7[yCIs���E����礻�K1�-c#Clc�.x��R#���.����h[�9�np%��p�l�� ��D&����MIbk�T	I���'	��[�A�
�qR�न&�-X�*Ī��f����,.���������s��O�߅$n�Y���ǋ�l9�B5���$�,cч�H*a�e�༂�l�W3L�1���f3V"�eaŀ���g:u�Ǌ�,�]��:�
b�©����`����i��f���2pT�e
�"��3_}5L;4�`�d��
+W���o]1�B�'"�D���+f\N�~N�T|3�lx��L�	e�/�]��BAñ��