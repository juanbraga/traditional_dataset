BZh91AY&SY��� �_�Px����߰����P�9� ��Kj&̔��&!��4LA������yChA�eѤ��� �     H�B�M=OS�Ԟ��P  @4 � �`�2��H��O�'�G�z���F�ѐ�  ��№nD�Sd"	!!� �@���Կ`%��QI�1#��C\�7�h@Tb�9�CAcW5�!��Eo�0K�ԡ�x��>O��������7徙�GY�r�SXڭj�Bh����=���\���$fW��ն�;��a��Ꜹ�r�38����$�Dw�囏���`�fL��s�~�'2��{���G��Z�5���F�0�3��H� �)t� 1��6m�]TX�؈�][~�� ���ֱ�RF����4�6wX��ZV$ì��seRش.��]]3Q�i�f�U�£��;�
�T�M�^}��n���)��������������Z��^Ռ�	Z�
�dRȠ��y8�.��1c�%\���6�V��TF���F^[��_K3x�m�j�U�$�R�[�k&�X]d%h�b�>�������1	A�q�'2Pm��U���QvK��Z�Гo�!��h=�2|6�.6�&a���&GєVg��s��l��c�t$�G36>/�W>��oY��8K���ƿ�������(���}�_�N{5�/u�=>VS	V�Z��-�:�|����Z��:���5�H9!	y�n�ɷ���&hm_�m(_��M�=�O))�D�i��|ǫN��ѭ%���)x��n�<����`���Ab��Je���860�~ ��H���XC�c�����^wL2�]Q�z_���Vb��x	�Bt��+8'���TdT�L��@8	4(K]��&��.(+������Ă���U)зw炝����$!*P��2KbuUh�!>M��G�
���*��qa��RѰ����}�̰��cy� �40̘lk��c�olǇ|$����X��@6�	w��ag�kf%�$0�Td�a��%��.��-Lh��I:'sHA�B��-��(�)!�&{!��A�,�,Y^S&�O2i���@�� ՛��m��hF�	r �Oa4�th"g���f� ��^�\�f^��I,Ƙ����6��*��k!���خ����!d2N��ر�8@�)R�V<vf�˖�Ҵ:�]��DM�$b�T5ǻi�ٸ��5΄�^آ�1U<h��j�a"%�j�%c'SQ�yz/d�j���[�a���5�J��:$�d��@����؟��n�鼖�E{��nN� J�dv��f��쩘�y@�h6�o���ܑN$)�C`@