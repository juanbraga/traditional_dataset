BZh91AY&SY-�� z_�Py����߰����P˛���E����	$�6�zCMM4�F� b�h4�&D�hѠ4    �$$A
zA��P��� dɦ�L����0Fh� 	��0S�(�=C�  �����-+ٱ$,
�$�!�\�$* {O�� 7|�ʚm�@&���d�l�IZ0ELm�6I�TՍi�}����$ss��0l
b,՘�T��f�9T���x�5�Z�Ȫ!�C�p��j���0�X�v��0��!C���Q��q�x4p��>�����!����.�Nt������/A`W��=a�#
�p�B�A�����w[h��m����=�X������ʝ5�1LZ����I~]	X�WI;��ߒ��/���6�: ��%�#YH�c�D9�B �z���,�jow��2t�ۊ���ƧbM�+��.�@�4$�{�!F�����Ű��i����PgbזF&_��UuNZ��H�0�-WS�10,N39u����N!X����L� ")�ep��PA���iqh�V�&���Sm:��j�>�X�d|:
���w�p�m���&6��82ߎ�[� ���V��Ƀ)�2d`���lb���Hi4�ƿ�(�lS��1N6ѪK�]�P/F��{���acT�X8�H�.e�vOs��I**��>[�Î������g�������İ櫮wm�~z���]���� ��*!(l���tb@jʜ�g��392��9a� ���^G)4��y����aF��j����
���X�4��"K{��D��񘲠;��
��֍���d��GQ`2H�2�JKϿjD��ce!���=��ħ����q�1v����|Xp3j�@�{���^U #!��4�(���-	�%P:�Fr��g� E!	+YxVZ���U���x��o]����ޠҚ�?���N\���4�
�3Ip�S����Ոg�w#�>z�Ţ�`�p�&`i��&��[@lހ�����HVn0̘l�g��`:�%=�)�f�r��`�`2� � ũu~��+]a�����+;%	I�M�T'�i�;䓡2v��R鐩���E҆��8��EֺF��X��Z�*a*�I�f¤���^[A><U�#q �
�:s�(aJC��.���v��և�F�f�V^�6����`�̑��l8O6���>s	�p�sQ³�p�P�D��(�d���0�-°� �P�($���ĄP�ӫt����I�wI)�D*�b��H��FI�\5R(����T0 �n�{`���轓�.)W�:fg�UM\�%Di9⑽y�/\��@~@�#=\wkq��q�3�\���(�ľ�t=���$ld��Ŋ���ܑN$�y5@