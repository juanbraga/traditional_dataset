BZh91AY&SY?��~ �_�Py����߰����P^qm�Np"��`I!dhe1����F�4h�&��z�ShD��=G��  ��  ��)�F���P4   42d�b`ɂd ф``$b���M�Q���ѓ�h�� dI �Ԑ*4"IJ��@����]�S;��$�X�Y����1!\1*����D�B�ڜy�cXBC�L��M ��*Bq|�>�^y�)Y��v��y��S���U�����#qZ�����iq�W_�VF�w��\I�	�,�����<}��g�b�Hf3b~���Ix�#a��E�3#���.��w*��z`��(�D��'���0�EI�u)F$�8V�Z�G.�VajL�EA�(�.��� L�[h.ᩙ]�X!�.��%����ןZn'̪�ufx��4HV��u]Sf��BMH~���6p,��]�_f��vk�3l� ނ���6���\(Ҡ�`�e"���ItK��0�	xU��&���R"0o2����l�U,���%]�(ǇM.%X�$33!Х��aF�d)(En��Q�)�B�5 N���g�d��`Q��( ڽ�$�c*�:]��Uj��<� >h7�>��;:U��;�c`�=A��������d.����Fl8���꼳�힛m\W�{᐀�MV�Sᖳ��8�Ts�%I#�`mr�l���cx��&C0�?����Tkm̘���9�{��q&\����9�l�s��﷨I�x��輰������D�s��~����X���D����l����i/+��2���p0��*�G���l����N�m-/)�D	�C�V~�T)�#rU�ߌ�%��J��/1�V�3��Q�k��)CY$�.$9B:e�y��z�)P�s��@�wIq�
��#J�݅7��x�$��V�c�XȞ��1R#�T����,r��� �9t�N@��Xq����ɮ�(��m3�J�ɤ��B�d,�iA[0�&�&t�J����(VI����bMT�( �
ý���՚�}H�$V����%Er����������e��6����fÓBU���<@l'�i�dp$�R�P�u�P�߰�*`��d+��޻õ����AÜ7/7�K����kH�S#�ST�4�Koj�	#���KBz*c2�ੌD�ɣ��c=��	���X�QR�������%�N�r)3X�ᚦe�dRM�w]I��jd�aj�~:���H�
���