BZh91AY&SYo�7 ߀py����߰����`z�]� � <z�YJ�JQ	"��OM)�=G��=z���1���"�P�P�2 h� �  U?5$�@�4 ���@ &����P�C!�z@=C&� �4��d�L����L� D	1Sz�<i5=<��z�2P�  ��y<�A�14QA�7!�,$��9?�xNdɐX@Rk>"xU��A��+!Ô=�&���F8o�,����X�4�4�%�%��4��T,,��Y5�#���Z�q���v�K��)����c��(g3�S.��dK��p�Phd�Ęb8JII����]*32�E�,k=K�\�X���CE`i��?�:�n@c�p͌�s9��n`�m���1��=H��65�=��lwwy���&FxzvqQʇ!��ctR�B�n�!o<]�Ot5����st�9�:���Ze5���S&g�%�����I��?>���E��D��i�ʞ4F̋�n^Bxq�8�j��6�3`�n5�5��`��-͉[-�gE
,��k�Y��56h�a��_�o�͗�5��6kX��!A�}#�хk-WD�a�z��5�y�i5����(���;|5Y&��b�PڝJF�x�  
ɚL��a$H��BH#%��)t.�����(�/.Į�����N�l:�hX8޸�{����)̓Z���t�ǀ��!C	�$Ė)t�]�x3={B�&%è��WT�ʕ�gN}{�;��dC��
S�Ώn���w��-�mY����M�M�v�n�=:�A�8n�ч0g��֢q�y�;\�?9daKs}²�^���HZI��	/G���L�ͻ��z}k{݁t��*4���mB4(k*�Q�oO�@֪�mCBu��6x��m7ggc�*vE���Gzgr��ŷ��+*B�����Jd��a�&�9QCF��^��.��E�������6S^�����m���/\&�}QECeA$ hL<��䶢�{|���o�d�O%Vc+Խ	���%R��E
��B��(9*$Œ��@I��aBD��G����V�ϩ�%���x4��� 6l&�kO%q7�f���LӚ����/��$�x��D�aH��ÿ��h���;���=B�d��ӳ	8��Q�(8�w��RF��ͳ��h��Lv���<E�l����w���i�:Z�g�X@�H2��
���Դb�$��'��C�E�<t�_�ƽ*9��c֟��~>���9a��t�U�V��R�)#ρ��Fԧu���ftʛ�J�V�_׈���`á�f�H�h7�F�a��P� �"��keCJ�P�|�$�D�GqS�I� SW7��0����
~%�uurb��Z�fK�t�A���_�����BN4�8�����L������ٸ5P;�4yM@Zm
���;ə��)ys�F���aN�ex�� Xga�0�Ո��>Y&���wR����:��v9�"�G�����惁��N���f��`�xQ%Z�C�wkv�H`��9
9���j¢�-���`�=��Ln�hĄT��:.��v"lޅbL�T(�4��2;�� JXL�˜ěnj������]�31\%qgU���s�<*2G{�V;�����`�Y21)�8���H��B �O2��(p=&���΄ �h��ȧe՚z#1`�aƑ[���GT	�[᠔R�B-q��k�3�*�Y�ƅo�U�#RՋh�����EQ ����6I�E㔘B����r��b�F��k"Bx�D&'B�D��p-�/�u���d��vp(�X�tj�١׾73#�ҥK~�5������������)�xI�