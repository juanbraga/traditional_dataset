BZh91AY&SY�X� -_�Py����߰����P�q���-Z@D!�2L)���~�LPڞ�!�mM��A�5?Jh@� h�  hj"�L���)�2�4OD4�LF8ɓM0�14`� Ѧ D�	5=i6�jy&M ��4z�P( �{�A`R�D$ /Md4$��V?�-�M��3�?D��q!�4�[S5����y��{�D��E�BZ�W'�O�Pn<|7�y֗�K����k7W�UU���b�����Ug��d����h�3׆3�3�Z�.s��˯��H�ؿ��(��������6w�$�Ub����ɏ����8��s0�<���U���H}��L@ �R������c�f�P���� M	7������qK�$ �!,���� �YUjh-��D�J��@�8u��fqoN��K��̳LO1���B|��l��D��D7��}x����,b�]�SMB��1�ڄ�!��v�������a�)�A�yNH!J�v���5�\��K6,�U�4s�z̞[K��2j�>���ի�\٦vU�j����C��TQ_�UI��ӓ�_!l=�i���Z���U�����fn&�?�d�"�+H�%�(XΒ��}ٓ�G6+M����l�9�w� �kX�O���Ư�YU)���Ƌ�<OC���-^��GK�e�A����qƟ	���i�=��y{,�Y��p%�y�w��R"5�m��+��%#@�I�@p���>� =�t�+	*k����ln86�M�P�
x��$/���b�F1�KʇQ���PhCGx�-�G��X����Q�'�7A��ݥ�A͕��[_e�)�=�՚\g�����^7yJQ&��8�����H�Z]��r͘��5���6L�f��hZ��ze`U�|˹��_J�v�PQ�#�Z{�2G]w�f�A!&�*����AG:Kf$�Q�Y�heP���4�P&bb;2�L����F�3�}�!r½y�y�I+�,3&��<yO�)���#]}ln9m3��j��$ۄ���u."��e�6���6�(���J�,NS
�,�C$��Q��a -#-zy7
�Ud��q�Oڡ\y��M�3F�5\K�P^�V�����2�����H��i���M\��ǣA"�%�,ſuA���<��a����E'0wmz?�@r���SQ�s�[�
���x�)�����B$T����=����3�02. 㸽I�R1��EB!�q��)�lj+��=Vm�,.%����5��
�D�e9	"�9���)����dM��n��a��vYR�lHO=����$��+��s�.JsҨ��9/5������d�[M��Z��s���d�7hW����w$S�	 +�� 