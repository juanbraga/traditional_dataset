BZh91AY&SY=*�� e�߀py���������`C��   wς�T�gh  ��W{� ���֊H֨P7���R�{�v�I�JK@j�s�wQU] e�-�4hcJ�1�Ӡ��Ul@QѪ��i ��=UU�6҄��$�TW�
    S̀�J�4       S���J���B14i�F�	� ����OF����`�i�b4 ѣ	�фO�J����4i�� ��&�$�$EyOQ�2  &�@ $�BhL@)�d�A&���hLOQ�&��OI��r�H"#���DGT0QUP�@Qց�{�ڤ�XADn�0=�����q�D� ���@?�¤����"7�V�"�8B�q��|�;�m�@����ⶡd�@
��H��VIP�,��,<!�Ē�$Y%abĀ�(
 �� �H���*H�
�� �HT��	�@P@RE�(Aaa+ ,`
H�E(B�
� � ,J�*�� X�H� *@���� ,�d�@��!XJ�*@��)& Vd�	ݔ�$����`5�/��B��Zb�M%�<Ѵ���y���.=��S�|D�]��U�]��ف<i6̆橕��U�MZs Q��� �]˱g'J2��B�TeU��3qU��56`dQ�Vd<!�Sj)R�Y.)�.)���y1F�)�0�M�(B(���хv�*I����r�&Q�ȸht�͋k�
��ӷk%��UN�K�ub�ӧX�X���8!���J���d�1Z��Yr.�r��V( ��sx���.,dR�L"�Ѻ6�Y�(��x����X�f�E���Ie��Y1V�U;�[��̄�2�.B��0d���!Rr"��� �����*�e1�`;�.�Ȁl�ںlf��A��;AU��B$LȺ��2�NL�uWP"�Vj�$D����Q�*��M^N
xZ��c(ؚ�A����J�,Fx�TC�F)�a�UM5b���E��E��3����q���dZq.b歚4����&�r]'S4��F"�U
2�\�����QI��)�X(O�X
�PVQaݫ��қ*�JW�A�n�*W�FX��vF�]YÔ�O�)ݑ3��SX���1��e\���	�e�l�b�F�"�_�NѶ�j���"��C!(�����rBs��b�ni��Rfh�6�LQ��Jfk왛�ff1Ӽe���M�\)Z�nӵu�D�A&/' �Ʈ�^|�R����͐q�>"0�d�e������j�g�1��I˼˦Qv�����6(K8��˼�
.K�7"��9��1�b����3�;y���N��`�H��tg�f٦\���y����O��\~�����{L5,8�9��J��n$a�i}>��7���i���w��k�����GYwaD�bֹ�r˔�E%ҺуD�U�@�:X��h��6��-ĺiw\��5�fa�[m��qͥ�x��P�Ia�TbsY��5S�F�])Ywh[kye���k+�Q�����c�*����f5�1����[cITzдM��Usk]�G��)0�)f�_;s��Wv�m�yV5�x�K1�T4�[\4�C7h�J�[L\J���X�%�2�L�"�XX�8�l�θok]DV]*靆�2L�yR�����-˶�`�4Ԥ[\�3eZ
�
��mssd�F
��tp:h�(�i��.��\T�;'j���Jr�2ԘYeK������%bC^pͪf\X�f��cU�#ݭH\S�C$˲��6��4IhR�j8�sP���R�j�������r����+��M��L�k��V�o;�(�*Z� �.�cf��X.M��V�&����t�z9�:zB,.� ��R�8�n�se����K�k T�Y\���+xM2X�mVܓկ���o�Qx�i�]�EՕ��(�k���^{3d��D���M�q5M��d��u�b���&��ۆ�����H� ��`tE�-��Yvʱ�5m�AG�B�h�z��cT���U��gIER۷�QXs���2����EX�-u��j�E��U[��ZZ�Nm�P��)�ܳ������TU�bT�l��:x��*����c�X"<8�PYX�4�P^2T���꘶��b�3����̲֬���VQ�m�pQ���L�J��a�C�+��+H��`�E�eI�Mf���-a��b�N%H)R�Y��R�÷����LJő�UTVQ��&B�,�TdS-F��fs'h;��T*J��U�d�R���k{�rŞZ���0�*�C]y�2�YV�9qB����2�T]aZјʝy�lP�dF��(��*�J��"ĝ҆��k/,��58��ͳoT��bk��9�c�*�����ה��a�ra��%?�?����DA@b�~�
��O	�Q�D枸p�/0�Ó���ƴ����d���"�ؽ�O���
�Po4��]-��+tIt#p��p3�iu�^Ҕ�mZ��a��X�(�j�n�7�Z��ˑԻn\�UK�l��,�Vh�R-��T��A�.Ԗ[B*ј	�
6�������� Ȣ$�$�(H"��� (@u	���S��-�g[��WMt��b�0�Ց��!����W�F�?d%����Xb�O�v�u���u7)=���m(N;�hu�CrXľ�D�uNv�\��<>θ��a�����`��mC\�a�.�_G�4VLq�D\n��Ym�*�1�7��x�Y�E�e6�5w�Eݕ���3 P8W.\ôbG���Z�*��Re`��6:H�8�n]}�2��0z)*:GPUj��w^k��*��b�Ll�NvU�5Vh�iSL��K�[.��5\^k�e� ���5W��s]�sXyO��uvC}�'�6.ǹ�������9�����Ȭ�1s?<V�^X��.*6N9�4[�����qUC�";B ���ѻ�f������}��t_:��)�շ"n��˗�|�o�Qa�9�����Rp��w#"��ᷙ{WF*������Ve4��ꣿ

�%^*P"헷�J���]V�gnM��n�٭�]���v�E&VVD�P�P4��p�n3�v�9х���X�3�q �o��{*
�/X�O݂����I��S�̳%����Iz�v��1�M�oC�����qU�t����7^mD.ђ��:sbM�%'�̚���<)���fu���y๝�x�ΩZ�W���Y��ʸ{N2�ʥu78,�\kux����w
%ޕW66j�&g$W�P2	Q��c��3�¨$�N'a�9a��*ڴi2Z�5�@��eA��V��N(lݪ�����M����;�apZ�n�GLC:Į�� x]=�S���_�;&|���z<1M�r��/q�]!�ΰd��� �\͊�Ύ�(���S
�0�RK���8~1��yK{8�{^�^V��ai���AI��`E�ɰ�5�&0���z���i5 �G�0𽾺a}/^>��~��O����j��W"�Ѧ2%��̲ky������xB(2$L�=9���l�ס֮ʂ����6	�k�t:r8�ʉ�F�Yɋ[�,e��	 �K0f�`"^gYQ�H�
OeF�\ʇ��L�=���q��-�����ٍ���w�f���=n�o �=Y}�`2�7ne�BL�`����l旋n�W�J�
�̪��!Þi���Y�K�Ξ���QCU �-��~�l�Lg�zUY�8��g�\h5kw�a���H�p/c�[8��:gLv����K=)����	��L�uԐ3[�\R�&�.�3���Ie�Eu���S06mbY[D9f���儑���ǩ����E���������҂p��=�����m_E�U��6�&�үh�Jv���/f��u��yP+�K`�0�E&x�-1���95w�Mv>{5V�qiTLƩϭ���Gh���e(F���y	%��BȪU�����WZ���'/ٞUƚy=�p	]�w$I�Dʻ�z=�r%��GBJ�,9�D�f��t��FLzj4��ENMu�7Y{���N2"}W�)� £��<�:�Q�� �O[���'EeE��l���b]39_V�i3q{�~v.o\AD�JJ�Av�]��y��Fn��UQs�ⴘۛ9,��5d�τ�B�����%�p�ưt��Re�^�5@�e�l�c5����[}G���S�3y�7/73s[�:�2]�8v��0��(Z�0C����m�����&�{J�6&�;�b��Mz���
�9OM�6�<2�ۙj�Z�̖lEe�c]E��Uǲ�dS��N�;�JUm//|2�m���u�ɷ�ǩS?U��=6�ar���Υ�\��dȵI���q�
�.�l^�Է=�sW��E�)K���=�|��M��=��pH���G��E�#�P&�L�M���+�7�kD�c�.Ā�On�~��= ���
���7��l�wF͌�/ӎm�g��r���=õ t}4�Ud#qm�-4~���Qw�� l����|k�[��9�x{���s&r�q���I�%u<�T��1�6�Tw��ʊ8�UՅ!	��-0���뗽Q��.*|+�ѐ�m�ʜ�iϬ�n�w1������:*�St��;�����Y��l�[�0�X��	�'��g�[{�&:[�1����C(�Fw�ꪥ0T�B��bf~Af�;�u�{F��9��+����~F�.���p���Ԝ�ryg�T�4�w�3;��;d��fsF��)�7���}�&�>����%0	n���y(��Vݚ@��qfe���E�IU�(�,"�5�=����E�5N��:��uO<^�a���A�����Un�������J��0�����5�.����q�yD���~q���g�U�i��M{�%2�7|	�d&�*��z�0UtL\�B�Yͅ7=v�=�b���*�Su�R1�5��s �P~�n�V3��l*�ܴ�O>	b˩v�n�������ߪ��O��h��
���dU�^1C�eTց��m��)R�U��eN�j3W��6>�{������,Q����������n��ά.����@� �������ޫ�V�UoW&{NƺA���f�#s��[a{n��a[w^�7ۛUn�.����a�q|�iW�O���'Tq��+6jD���Ú�FQ�4�L��=GJT��Xߊ8�z�ڞ��'ŀ��q��[3.M���pF��s}rlS��N�1j�q�M�Au�md�2T �`������ͺ�8�.x�_�涽�s}�b�ᅣ1�&XUݓO�᭟�U!�pSa^�5R���Eg��4c��Ⱥ�]�;�C镜{����UI���i���	'	3j���H=�f��׊��^�ʨCnt%7=ao���eU9�T_{&a����G� �)���e�(N��w;wA$���w:�f4;eo]�Г[z}0��+5��M �$�OĒ	u�W6����Rv�&�1�'X��MWVP���Z�[�J��vJ�ѪdF�(���K�y���q�r�]F�5RÛ�L2 `�	� Mڙ�V�_��eMz��P�v��n �Jm�Y���&���@zR��M���(j���[�:��=1�wgj�<�+@�~�J��#�˖��Jwm߂��`���Ud���������2��Zi+f��vn�뢳v�)�Ľ0��^mٵ#mNjw�M���u�)��eX^�l@���ԁq;�̥�#��]ƘՈ�bj�Fh���N�!�70r�J��/rhܳ7U�����WG��r3�f��2w�����TG��~?�  �O������ow��/k���#��w�f0Yl���[`;�JqM���t��^|�QW�8m�L�U_�j��RЄ���͉�nvj����Hȷ���*��\�˘$Şq��,6&�i5�T�2ͳz���n�40J�%�#��L��]��s���T�d�$��k��.�K�p�d��sR����ؗG�j�4k��!l�$ui����:^NN�^~S���l*�ɭj�5�5��es�\:�����+T;�������ڀ�c.1�\�jS�r9V3���ڋ����Ui!@�5:AQ����[����:��Q:�x�>7Rƽuf��T�R�i� �}���f7�q���{W�A;�J3��($φ�]�~i�D�3�����3Ttѡ�y��7]��ʜX�olVa-܃��P��	~9�?rٙ����ޣ\��;�.Dm�0�|��C7	{��AM򍼪�5��WOK51]�^A2�r�]���s�<΂@q]�f1��v�b�]y����i �M�yp�K�+��u�桯���E��"�Rk6���	�2\�P�z	�ʸ�9��Ӝ~ॊ"d�yE��!ub��ly���ɒ��!0��� }˩'��x��4 ^q�^��� ����.�EL��:Y�~^��5>=n��Q�zh���f�_����y�:)�4���*�E3�>��`i73L{z�����)%Y��V3�_��
�ψ��L��J�4��7�<���Fk�P{�L�=�ޭ��N��~��HHl2%��1h��x`OT���E~�t^6_E�T����kj�=�6���T���/T���,|ǠJ� �[�kTv2˖�V��L�h �d�a�_v]��^	^O���r����J����V@'WJ��Vj���{`$Cjj�`$ӹ�u�����}���0z�ٚ�$$Nmz�StR ���\�Z��GX�� vid���{�}�«t�-��p?3�G�#�AD�� #���	[f�a�"_k������C��z��=������:�T�νa0�q{/���nT+1a`S����72�r��M��i��8����n�B��;�77T�­T��v�A-�����>�!�8��Wo��$����ݽ5����ÂZ���Oy��4d�ߍw�-�'i=��BC�y�� ?Tf�.�����1,dɜ35��7�Y螺��W��Q�㚍L@	1��(����خ�N� K�{�u�:"XI&�E�Q����-A� �����B�w�.�J��H��;�����ڦ�ځ�6�״2u	���ߢ��8<3c}�Um�r2������y��B����;��U�Gd�㰩�/��
oKK���dNZP�^�R���[{q�Tde�f,q�$�364 8͋��;Q$U�or��Lŭ�y%QŬ������%��˵n���9�"�&֒	��'�m�,9�c�M�#�F��,^��̕]�4�ܩ�#[�.�d�~Țz�iB9��XΤ�E��[��.<UϦ}z��u��v#��#��W��f��ھmg{�(M��&�j#0RaP��I�&Hl�3����u2j)��i
���)��A���%��WG�ǀ����s_Of�=���s.Ȟ��:���׵��J�[m}q�"��q��I��ǅ�L�:,�4��p#ju6��	�r}g{ED���\.mmoi�N�t!.l��|�F���)�޹@E��ȹj�Su��e(F'f�h�*ۦ��1��\��雃�	����s&��\;N������k\#��
=ضӵOd�O;!�� )|�sN�C��Ě��{��`Ww�6.g�]7{��ފ^������(�!e��0¨f�Ȋ���j����+/,dۛ./!�C�v��,*�3u�Elݼ:�\y��'L]E�)�_O?��vJ�͉�)�Ŏs�k1���8�U�R��.ytM�PE�,"¶���CFd��x�]�����Ħ�8��G.�l(�d��"�YY��ź��٢�W��a�R���CO3E�M���))uF��R�mea��Ϊ׵{�1t�\��fH��/�F�1�ݻ\��C�[�C���dt��&�m����!T��*i]m.�I7]ZWDvN�L\����5�5�)wO��{[�_��2$֋�Ex�	�i��̼������tz����Q����3��$�d���t{F&7��Jl:o@Gzf�$�G�J�롼rL�K挥#��zd-]��r[�n�2[Z8���r�~D����^]�"�����e�'�Jpx�@oVEۚ�,`���K��Tu�A�/{�/��o���jE�]a A� �!L#P|{Ԛ�ar�6��x�9r�6u?0k�d�7Z�j��1 �̃]�4��d�rM�2���AI�^�b��wL�a!R>|�_�����SSv�zM�G�"�`Yc<���54����ʕH�z��G�֩=���D35"�.�w�N%W+%��yS�g�\��ݥ@Vf��n�:�bT�[w%ٍwK2)�S|6nL������q�s~5I
�_�O�Uh��"�zQ�B{��&�:%�C��g
76u礮�4��`�ҶIl��Eb�YV䉋,o�Lk��E+r�e�!vf\6 a�Qr��f�G������M�U<��t�M���@��5MÙ.��XᑤE2����9&���SSȰA���܇YUc_R��j�]&A��9�d	��v��O�Nmz��'>;	�N��3e��W���ಈ����n#��;^�΍I�(�-NZZkjfИ�-�z`�l%��(V	p�kh��!�H��y��	S�
�N�ٚC�6[xֈ73@*���>�����^v"Ꟍ{�w���\�:�j@�a^`��X�F�]\���e�|z�69��3�$��痜-Q���s��D7�Y�y��/ ͤWo���^����;��Y&Е7Y���
|����گ���O�(�W�臞����֊[%�̕6�.�E� � (I��j:-U�z^��5}+���׌0:�d�[���BsxL�U^�z]�[����6��{6c�TI�3�v�S���u͕�u�LN�>���`B5��� �2Uy��?)b�l����c1��q�ߟd�wC�:�z������;q7����i�
�x�Q�*�	��cc�M�ک٥�%Ռ�a�� �W�����Q���]Ch/�D K��˧�C�ǹ˪�Y|:����G���0zm����N	���esԪSlD�X�a�@���@9r�f�T����L�-��te�w�l�Y)-�Ke��;m����D�"�6�qɣz�w�(�M��m�z�W��.N���$^F�:�K~��mC��X�s��~�>���E�q��N�����C�х�����f�_Z��0�"`O��~�Ge�Yn���)R���3>R��;jkF�u����Y}9]����)�Md�[oFq�5�O�ͅ��m�����,��'$�h��lʹiʄK�EJ�+��b#�[6vX٘��UPYic�����f�aY~7(�Nb�C��^�W��F���KJ�h�pէ[�qsm�*��
���{�ǔ�Q�5`���Z�ڌ�4T�����dO����E�[N�,�YcLh((�6ͅ���1�*-ցe�36`���=�52g
31%�z�J�6�,D��"�ػ[f�/SU5K���l��ڕY�Z8��K�����Ǒ|S�Z�o��ۅ5m��	[a+I�t��n�L�6��y�c���h���x<q���4̀����c��6�C	v���J����H��
��E��W+��W�����8zw�1��U]ux�g'�k/�!���fv�ګ;e���~w�8�\�l6�ۑ��f�#�����yb���/9���cEy��9�|iߣ�8 Q`p�\
M�'�%���6�_fh�vޖ1zj;wۇ'�
�u\a��	�^��+Q)/O�g2T6���kV�6�H�4�_N޽x���b�b��(�}>̖X0@� ͭQ˖�=��1l٬�n""����+k����0[^�i[���y�5����
�^8��@A�l>��`�C�b�F����g6&��s�g����7�E��7�I��,�w� QAL���g_����lf֍�7���x�}F=;�y�$x��l��9��y�`8,��n�-��^�,��p.<��a�38&b�~,H1q�Q�e��ˮ2H阜6z�_w6�:�2k5��v���V�
A֡�����?�c\��Z�@8L��FHͨ��kZV'�Fpƈh6FJR8�Y��16�%I���%X�$l��S؜]���8�n%����W�ɌP��Sn�f5̦�>k�̥�D5��*]�藾s;\�������/��vd��؜�ى5�����q7t�q��T�[y"2D��6(�t�Ha�b*�9��4����g�q���8��?����Y���%Y�P�}YɌ� ǉc��T7Vo�-��n��1��Y�aP�wlV׏���	+:S<F�u�_��Q¨cOT�nջʥ�����.А���8��E-�*�.�5� 镏  ���`@h8$�Ts9�Q�L7��0z�f�_��tMG�g�y��CC)��X��UM�����zt�W7��˳"���7	����=oLN�A�&Y.숯E�����|zdw���]�YR�V���E�7
'&q���k]O���I-ǓM����357�3-�7�,�W:�ȴ_-�{��Cl�@�^d v��aF�k"��㑔�<�/@����}j��)��,�͞��f?�X���1�4X���]sC��H6��D&�	��s|}k��FE;��V��[�w<�x�Rը�Y����]2>VK��n.�˞�7Z�(d��ħGe$&��$,ӻ196�V��T��m��M�]��Kk��n�Tr���骘q�]x�1j]k��p��
� 0����˭���j�*~`�w]C��"�2�Q14X�gP �� y�w:�����i�8�r8�Գ8�;�u�d����w��<u���γ�y�}��!�hTQڋ"�$DD<j����x��0�z};[�1���6TQq�*�P�3-k��g�(��(ȃ%�E>J�� �ԊimY���TL*�P-j_�
���H*�_�
�a 8�Bj*IUF��#eH������:�aYm���ʓT\}aì�Ik�$�o�+�{L��O\���e? ~�P�w��?��qx�z�w����}:w���歉<I� �I�����4�wʜ]"a����;ί���,|kY�����~�GA��KT��"">�y��N@zr���/y� ު�?tH@A�-@�S��.��cW��S�8�͊����pϦ��v5��:ߐ��vٰG������<>�Н1!M�Kf��XV�f>���0Z�� ~�(��/Đ���kL��[���l��,S�9n<,CRIѿ6�Ԓ��H�V ���*�6�%0RA"�m@-"T�P�f�)B
*�PQ
F
 ���2�h� ��eF���B�������Z#�l5?�U@n4���B�Y699q�`j��q9������Y�;�I����d7s!�����_����ur0�� �ܹ��Y��mĘ�0?!3��S�����N���i}J��^s���[��:�/߬�V����N�]:y3�y�";X�D�zN���{nZޯ��j�>�vv�@�w�-@��;G�>C��D:Ny᚞��*�K&�o{Ĭ���(� q5qY@qqx�Ќ��I[�[Fa{�E Q���)��&|(q���X��l��):@�9�C�5�i�03��>jv��"4�	�֜��R}18ӐD{|� �����/�}��W�����ڙ����0lsY�-S����$+�DNR���<� dZDgF�!�ZPo���(Di��\2=�>�#X�'?e�k������B⮄KQ�ɰ��`�����t�7�3�G2:�L��$��l
�\�����7d��Z� �#��M�l-'%B�Cq�7@��aO��Ct�3D6r���K�Vf��;�m8�� U@�/Wj`� À?a��Cf&'�rUP���Y�蠿�}s*C�r�Z�w�Þ��P'i�ձ<������"�(H�Vz 