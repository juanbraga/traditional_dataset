BZh91AY&SY��E j�߀py���������`F�Ap   >    �  &p�
 �{���m���`*ւ�l`Z5)�Q!� �Fڊ�����R�E!�ZP-��i��jUiPA�F�F�EV���l�i��(>�   S�A3UU5 zA�2h���S���*S���@h �  Ji�4444L ��3*�B5L� A�������R �	� F��`  �&�@MS�h����i��4Q�&ӛ�5� *�C���*�� \�@h���I$�Q������!�������*0)"��)Y񸂨�5�@�ȁ�A�(�9D�����I�X<z�n�4E��JP��H�!t�z�F��
 䎑�
��
�i]�h�)#�t� hy!�B�)B� h]	@�t,� �PB��(H�H�x��
��i�i�:@�t� iB@�J Ҵ��Jд-:B�H���(B��N�4%4 RP+H=K�(��,A'�?�M�șxw@�ٽsT~�!�c�a�/ѷ�S��D$)qQl㺴��%�)I,�U�T�&��^Q��*,@�_\@�e1*�e� ��S0�&� �d�ff�f�K&�Q%1�?\�5Yfl}���4�-vS�UZ��b��PB���9YXe�RD��v&�}X�n�ni�y�Qa�3RѪ�n�dR����E��Ib��u��`����DDd�)Ɍ�ؕ8p5�X���J)چ�	��f�*��]M�N1�4L�M��F$�U��\����L[j��Ǆ��$ҋ���Wf�y.�㊬�&`8��}��3fk	�Q�$�N'�"2�!*���*��@�wV��J�
�W��:̓T⑓B�8�	u	��17B�e��H��L�Ǚ4��גE]ʻJ��Iݥ��4"�.���X�dV7"���R�ɛ8��L�˙l�W���Q��7c-�&�%��M�F1n�}� �X���#)ʅ�
j�&j�:�q6��E73"P8iM�X�Yb�7�ZOb\UKK�,g-ʁ����rXR��l@o	��WR��̹��E4D4#(���F�)�f�́x��2F,�2`:8�'2P1ҋ��4S�Z��)�3DX�U�nEa�u�UE�Q���hL;������5M�f]�m���Qt�N����UW�M��Ϩ8��D�2˷1W���BMT5uS��4��8�
%a�d�9�V���`��a)8�TfE�4ca�8&c�q�n��3>x��tB��RZ�rTө&UUT�;�a�(�I"C��-9'Q��"�J �e�J4�Ep�^�י2�s����� �B��2�z�c�	_�(�7l).D�s�9��Y\ˌ��O|����H�v���\�x��U���M�`]�5�gc%c����M5��\]��g��W��&�׵�V�l[�pbkj�j[�����]�-ZZE�h%-L8I�^4�x�T�q��]1ɘ�n[��ک��̣SR��Z�!�icYJj�8��ӃC-�ɂn�0�K��]�ݵԖ\Z0��UnMk�o-@s�)�ۍl.����mc�]u���ux��`��&��j�%��Q&ѳ$n��ͬ2����E�TjWd�˶n��^��Ѷ٬o4ņicsK��ؘ�F[H�Q�B�ΛKGhB���M�.�YV����W[�k,��j�Քً���;fS��pG[�@�hR�r�`���M���:�qu�Y,���Z]t�vL�h��mqF0+�mU.L7Xܖ�JB���as�n԰-�&�c��\�m.��X�ڐ�SL��kL�at��Y�q�;08K�È&Qfm�[v��Ƅ�s�p2ЬKYsR���a���t]b��ч:ٹ��3��+���QX,"�łE��̸�̡#�r��!p|����/ߒwIӾy>��mUQ�X�� �}����ţh_
�"d<y��Z�� 1�=\19�HUs�����&�﹍�E+��uukM�Լ��"�h��Z ������j�)-�ژ��)h�X���rNv��K@D��uU@�0���s�JM�Tw,B�1���k�����9)@SCBu�4�&�5	MR��i9:�k-��J5��]2�
%
SIlb\E/R��C�]=BR�iZ�h(ZR*��hCc4���N�EոX������:�T� ąT��N��%rE�i���]��4��RR�P4i4�it=O9���ѣU�����F�k����-u=�v�=�5Ck4���")�ؠ�b��՗��%W���w��"��
�}箽A�>0�|r��u���d<`r��>E���&����3�⛆e����
�Cf�C���1c�U��a�Kt�\���:nֹ6�)�Ue����in�b�
؅�:1��랺5�Ғ+Ԥe��0K�,6�04�uб�VE�Z��*�B�XPK�y��lCX�1��5%�z�f���b�d|NI!�#>�2s��{�|�-B�Sw�^`̥#�w^�Y�^��3��Y��9�f�)Y��䱙kK��-e^H�bie]!7BL��f&���o�^Y#�n'��u�����-ER��]ܥ��ۘ�;`2f��%��9)80EOQ�-�p�o�Qz~}�MB�*_Ajg�aL��9�b�Utf�o#A4��j8��ؾO��]jf�����%�'��P�j+.0�07(��!l�ـFY���b%�-"�������	"Cb{�nm��f@��j�ۨ<B��6�鉉�c��-K���4V�0%�"�s-�����v�eK�����E�2]�1�o"�u�Q3T"��������Q[�3.+%uP2�aev��ws"{�tR1�r�FgFM�� �jl�&dO�X	�!$��#��$���$�QmE�ۖ�ΫQ f�ף#mJݫ����B��"ފ'��
M��E%K"v���<&�٩��qpi"�*h\�(��N�Z"�����p�MXXQP������(P��&�_"�,#m�ٻ艜��Y4$�8C��^T�8�هb4/���\��VBQ4�� �w�lr<*�2�=4{�uE���Lt�م��s��;V9���e���`[�����(8�'ENbpjT-i�B`M心�������(^���:�m�j��#�?.�f����Z�^͝�'ed�ɨ����e�,�כy�F�ۚ7x���f�n^��n�f\K�Rj�m1-cg�Y��}c� �(A\����������i?�1?�p�,�R}�ꚕ^�bZjM]�D��Nz��F�fvv�>����16������:�\vV,��#ǧ��y���]ᛇ�5���E����K� Twz��W����4�ή癚*�-��W��*`��=o
��W[���d���h�lh�Ūc>�����=�>/�\xG�$!{�3��*&�4�;ڊ�4��Q�&��&*0�}�F��FYiA�*�œ�`MD��/��>D�R��~h�@� GnUEP��~�f-��٤DH:w^�ڄ+���P�c�,�Σ�L��6�l�>�b�]�3�����[v�~OYU����8�yCWq��o������.r�&f�y���LP�d�S$�A�E���U�֮�K��^L\�N߇��zA�|#��4}��S�4���X�4l(�����,y늎����j���а��^���� �9�Yu�d�ѫ��Q3%d��p~MAA!0a�/B��okG��4��Os��� �E;�0�q���ɭ�@��˵�-��V�קr�a���؜_=�SP`La�s2�&�pT���]l�ʭC���p����	%?�������p�QꞼ�SF�mϓI`����劗��\&����e��Μ��u^]沽-� H�����F��
��^n��$�TL�u�V]F9�&����P!ؕ�t���8�/E����
;*���j��6q{���5�탱c�X���{z�����1�a���*FA.o��sSF}-��}Rd�y��J���ߺ��Cf�����ta�s�������˕5�i%�*��Y��ȍz���*�F)8���!`Yy��òhne+��&h�h(oNmX�Xn�eU��1�[S�"�u����R"/�(���r�[m��l� meΦX�2b�$�H�#�ܶ�sn���FV乕��b�,{nn&΃S9�g�śBѲ��B�-4э��R�IK4�jK�,�+�F�1v˂&�/�Vy��o^��Igt���؞����y�d˱Z�JݙW2�Z]q����@#�|f�׿{���u�?aC��N���鬮���V�U�9�M=cs����Ϯ��l��H�|ȼ9m]���׎t� ��G �9���cr"�l=���6�
�����y�Lt]_�P�'	z+~g���קo�^�_zg5��*�~t'��v����:�\��"�`Z��N�֝�W�$?�!&Y�k4�H��D�����d����C�V�����3�y���")����]�D����qs(��Q����Q��!�W�A�c�Ld��=3�7�'
�h����&=z_U0q�8cGz�Vn��o�s��{� :@n`Ҕ",/[��Xhb���>0���2IEf���%�(���଑)=�i0u��ϫ�L�n���8ڒ�e\�NT�	�_�5��6<�/I`�6,D:fza��Ȝ��[Q(θ�wP�v�f��Ũ�u[w�f�ɓy���w���m�JS��p#;���;O[�u郂1E�IS�U�@[8��*����׻�_zo�M����S]T�5��L��b+ɤ�n�amLzY��]}��4Vc�D��ZV}�q�&��n��*J�PzV�
��N�x�����#�j86��w��:������z����S�,jJ5��j�i��)P@����Q+��g�°�	I�`%�]u k�UYn3@]���^��ySϲ���/BU["2�w2��A)�"yn�S������=�������t��b��?�A��y/����W��:�C�^����G�]�%�ND���Aw�>�S��~��Vk�JF,�$�۱� ��3���b�����eÚ���(3����]�8�I�,l�պ�b��)f�ɭ���r@y�2��V����5#5�6��n�&����'F�[uf'̺U��#"��aEU��׍Hy�R�E~G�茸>�$�=U?�Jd�V�~~����~���S�~�"��P�Y\��6HǨT���PsgM��^���M���V���aŃs�{xJN�~Ω�s�+!Ȫ7^�$��j��޺�F�2F|���k�������/`扼�ح����Y� 9���Є�R獋��h0ŷQbIJjke��bc5�m�
nP�Fwđx��%�^�bwG��"u���g#:�����cH���)x��ڷ�[G ��L����ieE�gK{s��k��Hp��oD�o��5�PO�lF�N�kj�`%��]�� ��A����>�qGJ�qg=k�[�p�A����:A^3iw��b��p졯vn��H�� dwE%1y�6��|u]:��7����b)M�~�+ݧ�+��e��z�h��=�غ���r�b`V���(�ǌ(,8.�ţ��py����^�u]*���ܳpA_�}~^8v�&��VI���:ﷁ�N�~,,��`y��A	6�a م[�l��D��m1:)P���pL�F��
� �5#�A�V�A
wEջ���<�O�e+��~گ��^�	H��'���;����c���4g��v�S�^i;����J�#���0���s��g&�r��2k*��sRG�f��j.x��w'�ƮK�
�me5����Jw�Q�W�oޝ�<x棤��#R����FK��5��F��o/�y�=�[���g�EdJ�O�f����[�ь.u�}~ޛIAL$��M����3Oҫ�c�sMs���N�s�F���DI���ʙ�ي�Cb�SM������"JD/�PY`|���o����K�3�rl�r��&��[�.7DP��N���L�#/-ʋ$�P��И�%�J��R79�,LZ��̋��Wx���q9j�qn�����Op�^���_�zw�o��β��=���6�=�W]5���^�Xۯ81���\4�Xˁ��*���:���^:��ҡP�"�nA��K6�� ��R#�+5�nܗ [���epʺ�Da����z�i��[�	)P�E�2�:[����kk��]�������6���җ$�ȮSj/r	���*�9���J��j:L;S�_8D�Z�g�6XP��Fw4T���a۠2||�U�=!�u�wf@R�@�`b�b���T�J��Gu��.�.F�ū0<�PP��vJ����b;�P���P�7�M����ݑ�<F����&��}���A�e�|�2��=2�[���3��[}�O'.��mlXP�Nݘ�I���AOL�u�]�="L;QY}�̠w�c}뎸���{4W�����}�"��ϟTR�D��0�k�Y1@M��/��ޛ��Ni6��3��4��Kn�p�6��	�m��_�1z�7&�Fqr����2�����/UJ�Tt�T�ǋ��K��	����#�'r�P�>Q�뢳��u�;15t#m0����Y�=���ӬA^A]�1L��V24E{�r���ۨq���gS�	$sض#�ص1���P\�S��q;^ds���ϓ��hT%��DW@z�m�.���iz�N�1�+жм�z��Ȫ c��y���%p�w��c%�4�V	#�m㜎����F �rF@K`�ݪW"�x;�ا|n���0��BG���̻�}���ȵ>�@�&t�<��hU��I������j3Xf��F�#L�$�����.O:gWE��)��}9S�9�ul�[�Z ��c�/nw�u؇k�Z�T-ҫXne��i��A��m��[6��TПN����.��>�G�\bu�0&���=�шq�c�{�Suo&t@%��D$�k�D��Y��{Ղ�����x��^�O�~��?q `����҉!B���D�a�uVˀL� �o?{������ʙO�IJ���A�r�A��C�:�j��E�)	˹{�4�A�*��!�n%w&�Ȝ3�2!��۫�SF���wu0�qF�-������DF�[��.���K���\;&�U`St9"�2O>��B���/$��Q��<&末��kg+{�z��L�ʮ|�w�wi1,͖�cG��E4c+%[�ᵵ�8�+�2��;��L�4_�s��wz�3t\�f�����0�qXc�*._l�\"mX�F?�0_(bM����.�ˣZm�u���R�b�����ҫ�]@A�U����kX\?L���lW��PIg�E	^�:	����un��p0./}�!d�Wz�1�uUNJ
VgR���I�.�}E\�H��ݣ\������˄�M��:pv���\���3��uRX�U	�2j����O�F觇P17N�ޖ�A��%�})�nJ������d�kue����cM�3P�qk[W�����;�h;s蛀*rc7�	t'�{��v!��]C�yp�.k�;@��>���Nƹ��n�ϺT��c� f4�xDЫ��-�0��e�$���z��	�Z���<��'_J�R�7�^�y"���nL�&:}q[������}�<���b�;z�d4��ޅ��[��>�o]V���+��
���L�j�9�������AnԒ{��*A�½��5{�ϋz������M��y
�D�&��fǳG.;u9�����{��ߖq:�d�t��`��##���=��%D�5U����J�);8|s�}N.%������v3��S$l"n`0qi
mo��Chu
�� "J=6�^���5�_��y귏�c�>��W���گ��S�m-?����2�U��7*�̧3�j0��峺�6�2^�GE�[�MN��/f�ٱ�	�[zgs')ج˥�0fl���!�n�o���d���ډ�;���ʹ�%�\��]����m���iez8�\YV,"Q���F�$+##4��:���E)[u���&a� �R3ivP��ajZ���K�(��lF���H�Z ��ŭ�c勔�y��V\@�k�v�xa6�L%Z�,�����&�:��g�p�a��&�Qڮ5�Tu�V\��V/b�r6�DI� �/�3�PQe���R�+��1�&�ar��v�E����2E�zcυ����̉=9>��7ؠ�=��җ#g�؆Dy(ԌJV�b�
�������dt��g�����D_�z�`]�1>kbi[���Q/=��%�a�=Y+�{[�雩3�v��u�I�ZI���VG�*x9`)�����:�'֠()i�1�w��3*�c���H��/�=���A������+{��֩�݋�O@[&-L�	0&���m��o6��I�1m�ư訑%H�H�&����g*r�˚��\@�����^UCj�Z8�j��w]�4޷���3?��%�9T9��7d���uGs)��7�o�b�Tyٯ3����vj�ч�s��'=q�xY��P
���0w�	�ٌ��D��2�ۯ ^��H���:� <�h���j�r�&u��G�t׸BM�?7F<ף'X�������^�n֩���r����uE߮,7�~���P��Jp����cy�6���=�2�/d�<��"���l�vx�Y��UA�Vo]]�72R�;��ێR�3>���zj��n_��e���uu�%��0�1Ԡ�s�� �h�J�9�NM(����	?��[GH�q�~���\9n�1>�\��e\��Zb�^9R�+1i�ާM�7;6��]�;3쵳�&<�)^=q���̒z�x�N;ڜ��S
g�9N�{����HmΡ 5+�8�����1��XTnIΚa�N�l��Ɋ4S��;NպK,��:*�Zlb�Є2�/M��p#n��������K����E�H2D�����5��6�����6� ��;=�s����gW�`�(ƞiP��rTy�&�ӎ3��`�2�s��m�&W|��'�Y\�C>p�N�	S���\ێ���̝�8�%U?K{�'��}�򨗐0E>���w��&��|=��e�`oj.��*���D ��%J�T��UA&N��@���=��5������?mm��]q�8r��^sڱPC��+ ���uܽN�ĺ�S�/{�+9�I�A��k��r�r�؞VO��ET����En��~���s��OMM-��wR0-N���軤���r�΢^���m��r��Wt�ʏh������
�R�r��~2���.�KY�v]<{ΞЯG^�Z�C���)f�bW-,��v3�σ�S�\��Q��9����mL��F�|���3��U7�`�"�(%Ն�-l�*�:�\
�6O���{���[5JK;&����u)�my���>�a��Q���Z������\K�ϖ��*a��Mf���]w��]�g��dVE�	Gݞ顂�x��Wg���,����1&N�0!�{�y0 �Y�n*�(��W�>���b������p��w���>�T�$�n$)�n��	K�0��gEcsN�E�f���Zw[9�G�pvߓ����Ęx.=�`s���|�T它�ɼ��W�ٸ/���ݓ�뗚��]�������iN6�ڬqF���)�I�=��v��I�HVJ��;�����^�E�,�x�u����R�$«t�4j�2��&���;�7��2�3!)��SXT�8L�K�6�Lsc
ݡqA��c]��:��Mqc���-Iuã�k�9,G��V�i�m;V�k5�њm��ť3K���[0GIn��5�#l�
흝���*$[v+m�v������z���&�ے^i��+�ҕIu�{cW���}��������ϡ��گǹ&�3���]u��h��	��}���\�͗eY���2ᠱ���|�mx.�E�oo�/[�]O��^��J�o_��Y[�S��س��u{�eH>󞻟rl�M�t�o.�۶�]�eӺ���U��u�7c�>��N����yS�,��'�X:�o�����ȸ�3~�H:�{�b`#!oV{q�f)�=�Ì
�0�=�P̞�'=}')���T�;}�+-�h}㕊����+?*QA3֩]]yVl���i�U���~��ԡy@�^����XUAݫ�͸���L�dn��JG�R`Ґx�[��L�"bg���m�']V�>���*�NU%в����>��u�wOX^�\]A��	�H��k~|�*�E���~RP�F؊ꨲ�3�Ezn�ׄt������¶%ۀAn*�ycr�r'�k0���̊=W	=��60x��ٙ幱�4j�gê0��:6�d}�����`�W�����ҏh��آ���nx,��K�t�qL�����9D�Z�|��:U�۪.��k���:R���n�K�&v%P�$��q7-�փ3nfrM�6�1
 $�p4S���cRU5��#��=��vy����eE<�{2=�7ߗ1i�XJ��rܮ��T��'�G$�����,�S�o'��n�.F� ���{��B(��oԱ,��1쒡9�+Yv�[���;L�1�N��.f2�&��+p�n��Lc1����m���0!v�B2bl^��j��jGiRTce�a��9UR�
�M���ح�˥}�.��{�	y�3�]��Sa��E\t��]��v��ڀ�-��u.$���3�X7�dY�x��6IJ�FGג1����
y��,A�&�C���{sև�4n<q3�H�m�E8e(I��(�јƴ.�хii��]�)��1Ў��W���ӊ/��bV��OWK��5�S�
�+M��"\ы�߹����ٳ�Ѷ'06@�+�G\wQS*�FT�Su���Jy.LUV�X6�:������Z�9You��MY�^c�W��V<�x����9�i2���}�Vxߟ�U
�^�W��	裎w�9�G9]o�я0���*�5^��a##&7���0��i
9�׫�K��������w������js�`̴�Z�e�,������f! 0��l6C^��1�>U�_�^�`e��\>�݅�b��iA�a$�yj��}fn�K=Q;ʬ}����t��j"m��6ñ��v�� �/�={�����&��o:�ǫr�_��{�^��&��9��1��YcԺ<&IYNb�H�`�-�v6�c*�u�3-U��e��|j�rcob�}��.Ī3�٨�y��O�j�z/aŬؘҔ�"�Ikp���ֱ�#�s�9�t����_����_P�=r���ʖ�� QQ��z�����?g�7�K��>of���n.H� �kJ�T-�W WP4H�@P�*�T��b
k��J�D���
����$�R�J�R�iR�b�TK��"
^*}�B���\F����@j
XFStP�!��1 :�>����M"��iY��1۶�p���j��5g�_� r�o,���>���"=~��
���\I`��c>�e	�`��L	���]
�A) �W�Q�ϕ1Љl͗�>G����,N�a��_�~�W���o!�>�X���Py�?w�ڇժ{���YG/�C�UP2H��"����A	)����<�5�� zӝ9apvE�u��͢�|������'h/ѷ�Q =�{�̝�H��B5�z�b��\i�p5�]�S�Ht��!�ŏ��Ԅא��Y�i�:�!���<uL�ӕ�^5#$�̺v�,�>�F�`@A$ V��P�
��`� s`�TTDT�)|�j�Xfb�#��̎��s1�kV�|��[��U%�I���M��~?QF��>�I"i�t�I�Ibs:�V���z�.i�M�I�N��
�=7-X���`>'��EG#&��Y�y�o�y&i��&���r!�z���ѷ(�[�h��v�y]���#�"��	��Hx���oNm:�;>}5q>eQ���IѲ[���'�0Z��+��Dצ��H	�xR<h* �;�EG�OX}i:Hzs�;�Xh�k&��J���"��(|�j�e À���������u�Dh|�r��2|r9�ybQ5�0�!��Z��S`�s7	%���Q�F�lY t��=�EF� ���;<颤�ポzEG��0��<'2|/������ߑ��~	�<OqG86U��J�y�'���>w���-/��=�{��/�*3�g���-)C�u=��%(��>�Y���{�`hy���1�ݖ�`�"`}�߄�̀�]����%���n~���d�Hi܎�Ϙ�ո��K��;�]f𬮐�r\;.�s6�ٶd�*7y��&���������#KsiN�7oݚ��a��z��k۬߁��Wy���ߺ,UT�b�����7ds��6R�_տQ�ҼJ���q[�E��T�L�O�u�z@�?������=$`�v����.�p�!��
�