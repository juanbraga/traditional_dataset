BZh91AY&SY6�TR �߀Py���������`�}�x	޼�iH$�4hڧ��1M=M�C� =C&�(�� �OMSj hd @   sL��Lф�hшd�� A)����hzOPP@ � �) Q�    4 =F�"Aɦ��zd#Ҟ��4yL�2 �ʩh�@ RdT	"�C~abE��zs��P� �6Ă�₼`�;Z������x}Z�M.�#@�W	J�Hm4��dn�!	��1��1���ÿ9LS�4��Z���gQ+JJ�]�H$Ap����tD��"IY�@��ps?#�N��%\�7���N����	�E��� ���BB	�9$�Z���p�-��*j6�:������0�Id���֬�I����F�/�wg�SR�3K9�-(���jQ"���&f���$w�a(EK"ڳ.`x@2q�q,�N�Q�U�����9͒�9�U�c)�h��c(b)�sX�'��U��i�geT�)�ҳP�T�qR;��,%u2RN�\}�Ĝ'��g�6絕�Ք�e���D�iP��j�6��/$����N��{�&����)��e��&��!����v%	�b�ٮ��ۂ/ ���+%�����Ww8b���(��ծͧ\������I+m�t� gާTd0��==��e#n)���J>ZP3�ˈ�.TXD7J�)X[[�K�[D�uC�\a�-�OMl��k�F�ĆpIUF�y�%ކʓٜ�<���ۿ/��q�BBKƩ TUP�[�XM��h�0\d��0�.�	1Uʊ�'EV!�Ɉ��
~�J�a�$0B��T�e�%W,(
!�8�zD�$ig��?tx�g�[e��0�� 섃���{�<�d�f�?ڲ��<x�Ò7«��{����l0��U ����i��&�P�ÜbI�7hsK�Tv�l�+q)�H�T�%,�8FٯZ�k��Ġ�������[�.�p�K���I+�&|~}�&l�-�"{��P��oS�R�,iQE�ل��[�l����NN�;�G��0�hV%"s!N�- �jW��^�O�����ŵT)�ܕ��5,K+v�`���(k��y.û����'�H�����g�D���.���a�e*�87�J#�v��Y�K^�E�<^��si�`$��6��\�fe�\�M������(I{A$z���X�\
����\=+���� P�:���aD@�%z��DP�)���Z��PP��qH��u���x3Vw1&ZS	�`�U�I���tg����SͬGY@8�v�#��-e;%����$l?�z/�5c c���׃���$P�{|��M�o9Va�$B�eSE��Ϻ���]��z"#~�HH'Ȥjά�d��Z��x:8Ȧ*'��L�<�U$P�C�$��������22K&@`�%�-ŷ\s[u�	`y��^��I43Fw������G)>�J��Va�q�¶e�Z�7�M,��d�8��E�w$S�	o�E 