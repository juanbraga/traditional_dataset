BZh91AY&SY���� �_�py����߰����`_W�����V���6�M*{djzQ⚞����A��dO@�i$���   4   i��ɂ0�#M1L� 4�S�I��z��d@�@6�9�FC&h�`�4h�2d`  �A	ꞔ�d�z�G����4ɣ"� j7!f�J
 �=�HP�ε�����H�I$��C�s���Af6���4k��}�Yy)�@�@HM�d!B !���b�}Z�z�a��x|8Lfj�uf�YЦG�1J �L$h��v��X�&���7�~�|kj�[�Y�F��q�+҄�BV4)��h�^��j�P���]��-���qI&�d�/��T���>n��/0��K	�X�펒&�50I�ЅY'\3�b"��;�U+,4�.0ᄴ�S	V�h $F���aF銲e��*�qX�GC�3��J�:�;��Q�v{����Ywʅ�)O�\\�yO
 (��n"� F�N�4v)�R�x5���ʢڕX�@�Zĉ��[�fv&�7�	L�!$��D$��D=�����.Ԝ^����IJ/W6Hb4"0Hl-�����5��%��*��-7�2��3����N���t:ѿ��Gu*�]�Ns�e�����Ōn�u}�=���X� A>��������Ȫ��=t�2_l;Y\�d�K��K�Ћ�Fg2�&��h�ij`���_Uj���|�3e����֜� 6f�OO�=_���e�g#G�g��_<Δ�5u�
�Gّ��7��E���Է�.�j=��{~uW��)��Ot�-��H��J�ƜU���9N�3�;� a�7qB�}�;A+�+�ZI%�҅������[v"�Oc��~ӭ޴lB��\?1���))S�!��O�u��	�X���Z=p���x���I�2�����$����ϻ����*(���9��7�K����t&8/���R+F�(P�u��d��\dʐS����f�� ���	4,'�t�A>Q�^du^�+L�i��@ʿ��6b&#~����  ����,�ԍ��v�jņWLw�h�Q@WXT#��Jb����f}!���gɫ���	$��40̘g����7<ǇL'>F15�Z���8$�I.n5�V�8��.���
C%=�	hP]&5U)�� {	N�
b� ��U�� u�J��No�GEPf,J�����MQK��Z��� uCv�ZltL̋�Iy o&�&�e�Kt��L;���:�.�}���l8:5��Ʈd����~	d��I��b�3�i�-���$�BO#��OU�.hZ��0�*�f���n�qj)�Q�?c�t�q��o�!Ú���V���-��X��maT�WF��]�;�j5��h��^��֦����w��L�(�o�}���Ž�x.Fe�+�d��4�as�lr�#��K#я��Qf6���ɐk�V��?��H�
8Y�