BZh91AY&SYFU�X �߀Px����߰����P�p� F:m�5iP$��F�e'�mL��jh4�#�bz�S�U        	
i='�=5<�4��4�=@  ��& �4d40	�10�!OQ��i�S��	��  4�� CB!hD�
2��E	F:�s�D�� Sj Axv�U�:�%f6��(�f\�8���}I:;d3����3;�����\�z�M4��a&$Q��H&��:�e7J5ٛ�<�L�
���p������}z��(�!+W�P�d��v~I���t���f3:��i_����ɽ����#?$R��UJ�ۙ���*�ً����q�!��d��Jn�ި��*n��H
6<@4��	"�)��1�$����)(�U9T�(�l�M�e	��N!��$�j�*�ELI`&��T[%�����'P�@��,ِ��X̊Ws9�M6%���\�.\���#)ZZÅ�K!!��tr�2(AD|��(��eE	e�h�{R����v����bIWs&�}�n"�J��$sR��8&�[*��/�{�R�2]i-�|�:���M�����H'���N�Gb�6+��2�m��	u�+��&;C"c?�\�_��1+�1! �cW'��\ʵf����rH�b��ٹݍ/I4������h�z�q�ov?-���儁!�y��r��IP���w��zq	3�|�_��(�L��j����f l��$�i~'��D͗���kt�D��$�|�sp���&��U���"�w/Q��:Ѐ�m�8��aA����
*�Ͱ	f�O�3k{��"x���Z�=f}�KO<À��pǪ�4�3�`��%�$��C<�r��`z�'�
�QԔ��v!����Y A|����_j�q���6Q,ٗ9G����b�/�TT��:!($�.��Y;�=�f��V�3�T���Q�By�����G����k]��^w&�hBvӤ2BZ��K(�*��U���U$�(*����\yJ���Bd��g�j�y\N*ZA�E6�jǄ�(�%������v�\�ƈ���b*I��RC�@�hG�G�3�fU�����<Zs@ްqJ N��k�AX���wC�Q]�6<�nS@k��gN;�fKAD�}���G��ڣ����A3Qa-� ���D"h鐾-ۆ&�2�C� Z0cKjf3%ᐃ��Ui< b��QLC���i�(�DT��	�0\ƪ9	�*VG#nGv�K2�3(��[��42ZY2WcX8d��.�p� ��v�