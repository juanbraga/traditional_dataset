BZh91AY&SY�uOu e�_�py���������`C���*��TH�>
�T�gh � w��w��[ (4��}h�MiE(�w׽J�邕�P*��*-�QΉ���U+�m`SF��4�#u#:
���]b�YR�1�@yk*KLB�lDl0��T   H ����ʥ��      )�@J�P���	�#0�144�2`A��UJ���i�i�4ɂh���� ��G���� ���  �HJj�������M0	�0`�a�	���&�M<���M#F&�6�MMf� �����DG( YEUB������|
RI* �7(�����87�0d> �#$��$�? ���CQi=�+����tM��;���ϐ�c + VY"�T!Y%@H�
�
 ��C,!�%B
H�J�
�!�@PI��I T�B	P*X��	���,��� P���V@X�"�d�P�H�(A`
@X��T	R@ �,�H
 T"�Ya@Y"� ,�X@B���T�P�RL@�"������|�hT����g[/ye���֖����D������~�Д�E��7��4��b&bmK	:�'(Ы�ud��
N�F�c.��<4̳�T�Vsw_'N�EN	9��Cvb��6��8�⑺�P�w�n�I3	d�b�"����-Wjr��(KO'+�eI[�n��b���Ҝ�H�Vq�a��*�کr�Q�t��pT':�S�в7!6a��[X򍸬1"^	6��A�U2)U	��Ph�N��&L��ه9������o(��5`����J������K���)�@�`�B�� �LEE�"M����*�[e�YwDe���c0��J/!��b��2b��.Ya�q*���%e`�n1�b��ʨ�f�Kv'&�^<�Q��b�6P��D��Դ#%����@�S�Ü��j�Eb3��W�1�f#P�/1F|��jX������ѫ�(w1"ܪ*��k*2H��T*YUl���`K��nҙ���4�ŀ�!erevm��拹4����"��@�ՃJ�����N��rK�8r�I�%;�&r�B�k�ݗ&1L��6�A1����R����\K���6��\�DU��R	��f+�BLN$���hX�� �C��C�4�*q�,�u�w��+�]-�����2��&��;WX�TJrb�r�j�]���0��)Jʋ�#�#f@jQ��k)&�*~�/��̺en���ʨ�b��3�����0���r(�C��s!a�l؛s,�%P��Á��?3.kY;kx9���x.>�z)䥛�y�~���%>0��יD�0���麻�����1;o��\�28"˸�
$��λ�\�p:)++�4JX�c��l���y�kn��K��uʌ[fe��,���^��K-UԖuF'5�CU:�jEҐ%�v����X;)6����R����ye[X�cƹƚ�b�,Qm�%Q�B�!3vMUͭw)ZĤ`�䥛F�x����m��^U�x�^&��d�(V�%���:Ҵ��*J���6l��*�VQ�"�XX�8�l�θo6戬�U�;�d����SJ��e��jR-�+��V��¶���F\��3Q��>�]��#J<Zu��b�Ѩu�HS�pV�˜t�CY�-I��T��I+1�S[��[�mS2��Ż5�s����jB�-"&]�4p���KB�[Qś��W6ڗ��T%�Ɩn�k����Y\�l�Je�X�f���x��͉D	R�1!u��5H��p�hn[��M�Á��Z�s�t�X]�+V��qX�`��.%���r�J�4 �F�0�]pV�d�Z6�,��'��4�����DA�K�Xܢ(��V��^�`{!(�j���N�.\6լ�&Sm8U5B�-�p���l14ƷW��m��ŤK �E�:"̖�i���b[kPQ�L�E<�,���(��lE�YĢ�m��V���2��%T�����5X��E���틻f��H��E1*��e�,�be�h)UE"�DX�([+4��v�V�U1q�Ags�m4����7�TQAv�R:�:r����b�_u۶ɼ�֬���VQ�M�pQ��C��J���v�HW4�+N!�׃�J@�Rs�NZ�2�ͦ+�T��+ٚL�.�:v�.�2bV,��B��iYD��*L5B�,�TdS-F��fo'H:�aU
���ª� m���TTCv�7�5�,��ul���W�4��T�M2��n�B����2�*.�V�f2�;u��7�ݪ�,r�ʢ����'T��C��eݘ���n�=���\��CN'7���Uĥl�]Ҳ�Q��d�9q�LJ{_���<�U"��|3�?����|!��Q�\�i�$nJ��n<�]���(�;ɬ�)�� "�ؽ�'O�񍰀��4��]-��+tIt#p��p3�iu�^Ҕ�mZ��0�լI�w5^7m��-Z\uq�Ux�έ�b��[,�Y���E��cj��H:�ZK-�h��VB�Yۘ`"��"�� �� �2�@P�(�&�뻓�\Kv�2�+��dp̱vɘ\j���B��?�"|��F=r}&�>�^8�VI��N�5a�ᮦ�Ce'���ͥ	�r��0(nK�܈�n��ԫ��1g������1��S��ӬAҍ�k�,6��k��2�Ɏ6h����-�v�]f<���b�"�K4@������򨻲���f`

�˘v�H�{��_E\]S�L����Im�K���T��E%GH�
�V 3���u�������h��j|˪�� $��%��K�[.��5\^k�e�Zz���� ܹ��9�<��@��!���c܌W�@�}PH��w��Erm�VW���+Q�,nn�'�-�cmeu8����U{gh�ԳZUWC�ɾ�Y�:/�u\��jۑ7ZEe���q7��(�ڜ�Y��l�8^ۻ��\�Tp�̽��x�݊BzL�	T�2�n��uQ߅h�(v�ۍ�x��.�m��&�F�Tl�®���;r��++"n(i�h|8A���K�f���ka�m��v(�aC���U��Q�|����Nd�ʤ�j���Y��ʈu���$�=_;P�ܦ�L���L��uL8�պcz�Q��6�h�Ss�9�&Ԓ��P̚����z/�gXw��}9wzA�@�����n���}6n�F\b�4n��;W��^b)7�j�w�U�͍���	���T�Tm�X�u��p�	 ���Ka~�R�+���"ߪ� T�)g:�"����]�^t�{�X}��ȁ��Ht����Ў�4�u�]!2@�{��U�迪vL��S��xb�f�֗��.�����Je���۱\߆����S�4��a���}/&p&�c����q�����;���6)80� ���6��$�X�/��CI�0�<������z��N+���|���3<=U��}��|��6�ێ��׹�/=���PdH��zsŇ�ى�C�+WeAR �wl�׾�t�q�D��.����|X��!LH�`���)	1�hp�,�<��O�-��75�E�X,�}~@k�~�l��V�;1��n�ۙ=��M��/�Cl^��̾�&;�&(�v��M��u蟏�f��*��3�ǔ����~=w��A�)��hx��DH,�����ӌ�z�\��3՜/�q�լ��^�#a���Ul�Ό�1�3J�,��'��ځ�a&B]u$��W�ɣ���n��$��#�����)�6�,���}�;�g������ˊ&����cwwyCߥ��{1%�1�ھ�
�=Y�I�Z�����խ�A�=�[�x�����o*l��j(l��(���s�P��)��g�f�j�n-*���4�3��+��>�J�т ,�^F�IF�wв*�z���80֡�����g��q��Om\��uݴZe���Rߛ�u�r"��IZE�1���ۼ�ɏMF�8h�ɮ���/v�])�DO����%4dG4�Gʺ*l%��mUC��²���M�L1.����c4����?�7� �s^�%w��v���È�#7E䪨��qZLm͜�t⚲pg��U�rr��t+a(V̙,�C1�%"���ƨ���f��v��o�|x��3y�7/73s[�:�2]�8v��0��(Z�0C����m�����a�n2�"�c�f͆[#|o���� ��NS��;�[��̹us-W+Ya�͈��ãLk��D[s�Q��>�S���awU�^��[g��`rm��q�T��{���C���[��?wc��Q��G(���\��b�ҭ���:��.j��h��)stg�O��)��G�z�	|���=Pi@��:K�i�to��C�ο5xqg�]NeؐI�m�O���raP}��F��J�3@R�g!��O2:{z���9�����:�!�l�i�����+�ř`f��4ϳ�^��n	�m�`�vf��ݎ��<��v{����n���clm���;-�q̫�"
�T�(>�b����j���|+�԰Ĥ�����}s�쐺�ǞWm�@��c��U7J	���j�ڼ��o��aU��	��@��z���}ŷ��c�e�����R�!�U�xNӪ��`�S�q
*Q������m�y���D���z�S;���eػ�Ka�&��Rncx8�\��*�~�=���ZJ3�6==�x�fߥ�=��s��^��@��$9���%��m[vi�řqu�]7����:k�ʳ^��۶�ة�^!�U���Ղl7@80>4Z���]��Ë��6��9AR�=1�3��U���kޖ:ۥ�.7��Xb[�̲��(�/hwr8eln���M�UY��� `�蘹<��+=>v��;���(_nU-�۬�0�k���4A(���~��"�g(7��U�i�|ŗR����US-GoD6;<��D�p�ЁS��l����(z�⪚�>���q%*Z�<̩���Fj���կr^9���64���t�r�^��^¹Ձ������=�E����D%�+�꾪��iu{kz��Z��ӡ3-9����p�E�k
ۺ�Y���U���m����r���V�����x���1IVi�o����at����k�(npa����}�,o�Q=imOV_���zĸ�-�� ����8#}�9����v{��C�-[�n5��sH.,ІJp�%B&H���<�۬�"�e��kk۷7��+nZ3�a ��]�4�����Q��W6���d��T88{�g�#�QS��2n�׻q�>��:eg�z2��Rj��0Cb�/BI�Lڣ={Rp������׳r�	���ol���=�T��=��Ǹ�_�� e0cr3,�E	дN�n�"Ô�kV���"hj�ڪ�>�Q���
�,���#��ʪ�CRH�f�4��uH�Jp���\��a���.�Ī{ml��չԪgd���Dm�`���[��wOW7-����`��U,9�TA0�p�&T87jg�xEZ�~��5�71B��m)��%fk� �Q�u{� �)D�&���Â�5^lTmW*O���H��&j�9FW��]MT��hG 3-��A�v��!���H0j�d��ᕳo<������"��+f��vn�뢳v�)�Ľ0�k�=v�����p�7�?F�~D�U�ۗ	�R��`\?yKdť}F���O�9z3���:*p�k��c`�:�J��/rhܳ7U�����WG��r3�f��2w�����TG�����C��v~����9���Ͽ�h��>�g�~
9��/9�j2�1U�����,WM@/E��q!�ӆ���eU�`樌�-Km�ؙv�f�ͮ�FE��t8�`AU\b��˘6���n�S���êGfٽnqƋb7Y�%\Ic H�S0h�hf��,�A�e``��F
M	�ɸG2jj9�np��T�K��5Z5�搶W�:��e����NOHI�N���g�aT�Z֭cZ�X˦W9�élLҵ@��}<Q����uj�I�w#�O��D����5�[��䑋n��� ��e��Qp�\j=�R=���S�m�MB�}Ա�]D���>��f�5_`�;ٍ�\@�37��ŐN�p���w
�3�_�{�4L�f�z:��4h`^A�W[�q�vv;�^��J7x��f2*{���撻O�}g�\=�5�9����N�y���7�囍������x��QSR��mk֦�V�OT�y3��?Wj�N���N��v�#vN���6���=�C�2%�HwC���`ۺ���?2$0;m�J(��I�ڣHD,1�	�2\�P�z	�ʸ�9��Ӝ~ॊ"d�yE��!ub��ly���ɒ��!0��� }˩'��x��4 ^t�}'-n 'L�`�j�E6��5��|{ˋ�Ӷ�2�@����G��M1{5[1J�|tS�h3�nU*�g�}W���m�C����6��b��k<�d��;|����\��m$�i4��A��:�cp�#��z�3��D��6"w}�^�p���&]k=�\be���b�I����)m0�IG�·^�0`�V2�{��Mlo��v�V�q�|�GS��4#�����I5�{mj��Yr���I�) �%��{����uR�J�}D����ϊP�v�j� �:�V�:�P`�����"��V	8�{�n�W��	�j��ݙ�"BD�ׯ�7E  �Ѭ�Υ�=u��f�J>~׼)s}����T\Z�����A�c�D��?��=���0�J�7c�}=t�Wv���/���dL����0�ݏ��ꡑk±)s~bs+cܨVb����:1�9�ne�.噪�3�)�(�g�qk˜ݤ"���&wrnn�)�Z��Z��[����G�YQJYo�E$����ݽ5����(�8%�����w�@~3FL���z��ڒv��hT$>j/7av@��e�Ó8{3��:T�Y�䷎t=��3'��G�k��jb �I�^�E4��f�v�w��������T��lXe���D�Pv�<�n��z4.�,�����32w)w�׵M��~m�hd�0%㋿EY�pxf��-"���b�e�;y#���Vo��,>��Y n�eU�Θ8�������}G��×dNZP�^�R���[{q�Tde�f,q�$�364 �wpgj$�Ą��ܫ��1ko^GITqk/�9Ά:D	`8��[�(�w�I�u��n;g@���b�z���G��ـX�5Q��<��M>w*z����p�(_�&��%P�f��3�'�f���v5&�7��^�L�����B8Xi�;�'ܼ+��#m>EF!�K�8tF` ��f����M���3����u2j)��i
���)��A���%��WG�ǀ����s_=�5;�'�lv�8{�k�~��{c�O��r�g�n/�5�YYB� w��) ��8�郖�E��F�nb�N��4`�'=��}�/��R��n����
x�;<X&|�m-VǴ�(��-*Mȶ����[J�t��p|_��~��Mm�����VD��G]`MQ��g#Ӱ�d�X G�bϙnl�O�F{��)�3<���=���c+B��$@���]�"��8z��U�����G��ޭ��ފ^������(�!e��0¨f�Ȋ���j����+/,dۛ./!�C�v��,*�3u�Elݼ:�\y��'7n�~ӿh�<��0;%L76&(�tK3���lF���v��7�]q�j����]iR��6CFd��x�]�����Ħ�8��G.�l(	b��kRcdl�7,K[�c6�w1]4��Ӝ�S��ܳ�ޝ�o}��Pѵm���[[)i����
m��H��s�"N���z����f:۷k�Cc��y+zh}|7^�j/�&RF����joˤw�m�\۳5�Z�F����ɋ�Y<a�ƺ��E.���ku��t�D��|�� Y:�0z�����rջ��c΁�Q^���7 u���=� �8z|�щ��|jR��ǎ��ޙ�	9��R�z�o�9MN����O�����k�X�{�fSQ�<�u爹@�D���쌭�g�.����*��堖����@��E�u�����=/�{�!P=�z ���H"~O3Yԋ��� K��^��	D-��(�� t�}'��I����,��
.~-yn�t�ٴbA��=id5���Te�9y����ެQ��靬$*Gϛ��}�"cjjb���I���d]��,g�u[��+>��v��u3�Ss�]_��	��^؅.��˼;��	�g?7�i��% T�b�YV���vݓ��<�����K��dS���lܙ=�{;����"j4I}|��ʯ�R)W35D=߂i�C�A�7<����Wz<�H�\{��;8k<O��6��0̲E�!JܷYr]��(�O#��<T�p���}^�ɽ��=�W^]6WϠ��©ĩn,��k݀�*�j8��q@IU�ͮt��0+���;*��{����@�kL���^zS���ݗq��g6�f}���'x	M������G�����YGgO���3��{�:5'�$�9ii���Bb̴2a�5��VءX%Ú������m n�LU��%N�+h;;fh$�m�Z L�`� ���=�}Q�w�".Ҽ�E�?�J�Q��u8ԁ�¼�m����������X���_-[�m����{��e�5,�{<��C~��'�2��Ev���U�n����ٳ�l�]�{:�F��KK�uuAmW��Q'Ôp�z8+��	�Y�%���I�$�i`l��j:-U�z^��5}+���׌06�c�k��;ɗ"���D�L�Τ�I�\z���y��T�p���D�8r�uͿ�nl�5�>���`B5��� ����y�����K:�\*A��V�S�V8l���r]�UPt{86�n&�����#�����W��~�Rr��������S���:�RS�޼C�֙��;#rk���Ư�a��t6���곫/N�{{�:��=�����qc��+d�O6uE�.�
������Hw�`s09�����7b7XX�P�Iv3z���oT�{͘k%%�	l�y��y=콑'�ȮM�rh޻���;�s�G�h���?K��%=	�����߂;;D�P�\4*��%���z�w�J�ʢ�h[��
�!wFK��afsz/�ݪcV;�6T��ht��=��e��,�J_�bt��J���9�H cp
F��9����T{���y�j��ޱJ{5b>���lb�T��(��Q�d�1K���R#2�br��uȩC�Aeu=�Dw+c���3xJ@奏��g��ݛ��e�ܣ�9�5�{��^;y"�-*u� m�V�nE�Ͷ\��{�*�s!�C7R�EFdՃPj�)k'j2��Rr�N8SP�B�Xn,��9`��b�a���k��ͅ���1�*m[@���4u�Zm
uW��	��3�����Q�U{"\ؑIl]���ۅ�n�q]R7M��R�h��4�0���<��<���9iC��que����m������J�}8fBPO������>�,!����c���6KS��;��� )��bT)_l�M=��m"���Qe���.���c��̜�~�̊WW[_9���o���c7~�����PF.W�TV��	!>�8e�n�r��Q��w�ܼ�]��Y�_f�/��Ɲ�=ӂ����[�|bY�*�kU��U�f���ޯ(��}��q�*qp�gU�ꠜe�@ҵ���vs'�71�9�q�[��*��u};z+�Y<6,F+i1r���z��ָ9��i�6-�����() �0�.�SD���N�5[]<��Æ��b{���3�䪵�S`ƱF{z
Am(�S:�.���߱��{=��۾�;��Xo6�gxo��AI�![ـ�[����&��'��^���
oY;��9N��zw�H�5?ك�r�3��H�pY����[���Y[��\(YIx� �>m�no���	3+|�#��i���:ܼV��0f^_H��e�o�I4"}�d��0	�XM6���e��-���ܽ7%�=X:,�p���0���F����<*<��`�k'ޕ�庈sh�P$�z�r5��ǚ��a�^������KR���e`�ٜjf0��;�gnd[}������ϟsB<��M��+�{(8g*��XZA�fM�͉ȝ��CQ��z�hݧwJ��H��#$NP��a2���HԆ�6"���SOlmmf}�b��k�3�!]n��c��Kެ�~DA@Jr���\,��6�گ>\Vs.6����K�~�R��ح���Vt�x��޾3\@��*��=R{v�B̪�O�]ǽڽ�=6v� � ��t٭�L�xi
�Ƭ�T ��fOTj���b.�/0uW�L_r��u)�)�-�X�}���P�E;Qr(y
�WG+;��.�<�ږ��'��^8��51;� �d��"�VzaÛ����]�Gv+)�Ы&��	��n<o�)>T��p��#5����D������;���7��q����97�eŧb��j�fy87� ��p�Q�ȱ<x�e:�=��!`3�lZ�3�n�3�g��Y��23^1��(J�'��'0�Ɂ�5�-$�e���!@��Kg���c"���+�6n��M�8�q'��rǰ�;u<neBA%x����4j(c�^凟��wx��Y�3�r��w��}@i�I)*��mܓ��P�E�9]V\t�L8���}�.���8
��a�uk|n�:�Y��Ʈ§�7qU�:�2(�\�3NVu&�����{���W�(��p?2�q��R�nn�����d�VL�Ô�Qtv_�~���A�z����r�Q@a��UP�^���R����Y{vW���"�+v��aX6�,*)|L�|`�@Ȃ�l) (�����pd!�+)!��L�I���%"���*H�!X�T����I(d�CI*��K*E�숭��] 9S�ja���C
&Qo�����"�*�&�&������S���oի���U=�����{�|��2����_�_��G��{����i��zvw翿�⮉<�������j���j���W�_��;?U���35���������m>�Od�p���`��[��P�g��+���8��9T�C0�$  ��HJ?/b�n;�4���Nt��o_h==[��4���~c�k��}h ��ؾHuNt�\i�
5���[4}{5
X+�& ���ҥOQ~i���L��epoݏl4��퉍+�KH_
$��,�)*�>�F�.dT�� �`"�� V�#Ai@���
�A�PX�X��*�"#l.�T(�(e�wJQ�:�a��Y���T�@�+@�Mn4`d8x6��BB&_w-1�(M�a~����9��\�Xut�S�ԥ.����� ��\���W{F���/N �DǓ�K���m�2k�����<�p<E��y?�\x�/ݙ6טޫ��˟ៗ,w� A�q��Iɜ�i��	=ו����e�j�Rz!�7����F�P ��G�}o������;)J�(Y3f��JXJ�@<�eT��xV��SB˩��X�Pq��2&������e�@O�����v	��[�d�Dс03�q r� ������'Jt��B��}����_7a�܅�-�϶��}?<���&'q����foJ�t�~2@�y��Q;N���aFs��;��e ;NXn	@A�����1��f%�7U�h�ɐ6.HB�.B%hx�5�6!(J�)Y���Ί��]H�G>�g���u\9�Y!v���d݀^��\�Dl�h�ڜ�%R�CD���;Lzfi3���x��M�)TկQ��ԅG�M��l*�ы�ܖN��w >�]y��v�*���4���@��vs
!��ˆP���p��qJw��=i��_�]��BB=�=�