BZh91AY&SY��B 5߁px����߰����  P]��gv�KA$��4��4i<!0�4�S@i��i���Bi�B���z�SM     �&��B4���SC#A�@���L�1�2`� 4a���)�L�d��5Q�zM d4 ښ5�
4"BH*
���[�~�4��;C]��n�0W�mF���Uz�-��5�3�1�c��虫+�6�	�����C=���q%��؜c�$J8��ac;x �,�%$,S��E��֞KM�9.�i���<�*[�p��T��l���h��1�96�3��Y`X=C52��A4�;�(,k$�ReNԵd�e�"�>���Mi!!%�I$
�����0~��.QS��n�.+�˚ن
X�!�or�6˨:\U�� ���6�a�Clbv����d�%�i��Źk��y�Qe}���t=��󄜒F9f~mz�rMb�}zx^�ĩ��Y���d%��r��cgLeA�-�qX�%kN��?0G}ǐ�B��-��^8Ӭ��&��B������fһFHK��8���b��P\0�W���cmb`�dƻ-o�*!�)��Cn�}Lr�n9~�[yuEK�Bp��ɖ:�;*���4�&��i���B��a�Ҡ�Y��я�.��r5�>s=��X��00��+�թ��ХG�"��e�7�~�˗9��ZMd�b3�������nh�7�.�J�1S�7b��f��h��fj����M��W���j�ɩ��Ì"��C��S�DU�1&d/��I&N�p�#�����1�����C&�T\��(���.QǦ��L��
�&?�+٣�:f|װ'
m�8��3���1�rX��gɖ!-	���s�.�r�5�����=�J��*
@F���L������̢����s�
4\*"嚗��t���f�mE�ehV�JTN����gB��7�U���20�R[�yŅnWO�^�N�r(+��?;2�T���LƦA�� ���	�|����)��n: