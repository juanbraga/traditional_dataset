BZh91AY&SY��� _�py����߰����`~x�׷D�����jv5��a$���1 ����ɐ4�hai��M&I=)� dh�     9�FC&h�`�4h�2d`  ��)�)�I�( 4� &�   E$A4�CA�=!��@ h 4��$D)���oTzG�=#F�h�  'P
� S�I�A�U$�Č�����(e�L3��HfJ���tI�ʆ�n�ϯǝ�0)��I�ӻ����`cu73���[E�z�uk�efz�8�K��[��;��p"�Bf�D���\��?�2n���fC�m��
������e�a!�di�����D��iBH�����m��hg8HV�0��r��Ґ�$�����6gv�h����6�]a��!�(:�wO,�(�~6���E;��T��f��z��0*ːf g��
�`�lrP]ŭ:5��!�	sk�1"���wu�^p�b��C
*kF|��0
�D�y7�����ƚj����]b���D��y �w�w� p�7Z5o���}y�O�)�S�SX�ƞp��ZU��K*\;  bm�b��Km���A��u��_
���m��o��T�ɐ��[���i�B�C�����lU���׫�ČL>&
��^�1��}�z���c*�q��^�*���uA�&w�'�o"#���O�U�q?\{R�\@ @r����S�gqN�X&wF�ULՙ|Qs��R] ���ͱ�.j��Fڍ�@�����$�1`$�U`��'*�)%.Q�ɷ�*  �'C�־z���;�xj�-� ��t:��{���9�
�n~���uF�w�G"���>=�[��Լ��sY���)��I�x��q!���  �f�ʀ⡾�`��^��
P�
�A I�|k�Q>��f��Y��LS� �q�CQ� ����q#�U�ҙ��;PӖ2u(��d�r��B厅ϱ�{�+Bq�,tcZb�<�ӻ6��8�:tһ&Ô�'vaU�K7Ƅ�kJ ��[�S���-�;F��e$	�%�Ιqd��#qq���s�Uʝ�N^&ܵgK��.�oÁ����5���)�������GNKԊ��)wh"Zd�[�Ag0;j�0��2Y
�T�W�0̘k)�t�O+Sq�9���'�c9�J�f7�#UU�u��$�1AQ�lJp�A2S>&!��v��S@� {��UB����j}���U(3�!�6?T"D`+�VgV��
H@M�K:�29U���'-�Hl�g1"Ԓ\~�tx0�,��0�g�U�~�yn4���R�DC�w�P�lZX��Al޴�	��V-V���!��Zh��)$�i�9��Q������)�jX8��3�V��'�Q�翁\��`HE��T\bU�W�Bp4�e��,���6���sw�#P�VÂk�*(U�"����$LC��o��Y�j���^�c��JK���-�]_fF�yW3.����F�q$�cLF�x����.�p�!�3�6