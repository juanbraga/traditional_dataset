BZh91AY&SY9� �_�Px����߰����`�&� 9��H��T@�$�d�с&D��<�!���@�� ��       T�0j2`���b��ɠ�`	L��� 4 � s F	�0M`�L$H�УjmSz'�<P�=@z�'�Sz�HBF[A$Q�@�I$��Z���(�ʴ��HCPÉ�YAV6��M�h*�us��W� 74 ��B[3�u�sS�ֺ.�$�����i�$��	�N�iT�6��T��GAKvTR&�ۣ�Tr��a�\��H�J�c!G��˦F�t7J��p���! �t�BJ���=5]�O�HCc���N�?{�v�i��0�'��/��#���\a4���$�r�=Ԣ��UZ1�m*%	G;,�4����I�Ĉj�J.B,ՙ�b�)�S�Cc�wA�ɤ&����i1����q�+b���R@|��P���WZ*��6�uT`I�Y����YT�ܕ�/��H���N����(������P�P	�,&��0fr�AXӎ�Ll\,�$�1��U�������=#�ŭf$�-L�ҥ%a陗 �Id`F�K!��ZU"�C���Ԓ���D����ǔ{b�y�N��g7E�����
��}�,lM��l��]>�Y�)H�arU�&�#�Z���[�Ԑ����HD&"p��'L��׊��U7��D�i�Eu�����䖆�D�c���0`��~�Vch4DT���1Z#�ql�.�0��v�~� H�.��"��
w�D����hH�3���-N��$��=M=�L"��xg��ݍ�!�~s�Ezlz�||iBc������e-1�t�h@rT���Pk����f�Iv��F�ĄyCiB��A���4�iK�x)�p�_��R�UrK�P��w�����|�^͈���`�7%��B(1f#�{Su�
y�����]�l4��V^�C 窙����sD0�G(�!���Lde8'�¨:d��"�� ���.��^�&�V]����f)�n,J/� B1��5#��m��Q�7�$"�7�ImP��7�im�ᲄE�'�e�:k�NT["�IQ��Mrȩ�nx�9D!<�m1��Y�>|����S��su�A�6�!\�x�:-ci�s��4�"��P��h�jd�1��$�L� RJ�O�D��Q(-�jI�3����.�%�QVI��@J�$͎�qPHD"��1��GbMX�QX�����bK~ڈ�����M҇���|�蘳�� �.�GV0s�F�a�:���X�������:�I�:N���*q!����K~I�0�s2U�4�z����Q=��R���oI��m���_ie�Ʉ��=�����`�tNƬʦ7sfC���43!�<��Yg�6���ٖN�!=8�q:0����e�������F�Z�
�EԚlu�"����Z����V_c���L��-G�]��B@L�W�