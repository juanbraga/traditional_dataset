BZh91AY&SY(�g� "_�Py����߰����`_�ݏN� ��T$)S�(B���zI��&���0���4i��=�5)"�       ���� �A���hh@d�4@4�4444  �  3�##�@d�i����2b`�$D�hJ~�<I�?I��D�4��#@=C��5PHV�hD�(HX?���%	��^	|�;�bGz@/k��N�$ 1�X�=L���Yg����ז�:7L�r9� �
	������DD� D�  RT$�H�F}L�����3̟e����6����"z�ߛ
 �W$lL �UM�ZVR0�N�]L�B�J2p�4��DD@�SyBr�P�P	r�u�{dc|�</���+�8A#|��֝}ibQ�J u�I��0�0;��C����y>7��|V�z�m���[m�m���n�ffe���6[m�{�������{��[m����wkwW��G��#�� U[Jrm����c�h���[��46��o�:9x���͋s3b]v�$�MY2}Ǔ�!��x�B��2�@5�v2MC���b5/Z�)K��Ի�Y�C�'mĉD���Ո���\��z�&Hq�nG5�)X@Qh��� Tp��׼:�\�����z�o�$�M�]�# rub:�D@F+U�I:@�pî�Z�NRR���$mI$�I'Aae�tx'S��5\؀+*L�#w�hƠ�W=ѕY r/�
�� �����^"I$�&�M���#;!�� O��=s� �!��.��]d��p�[E��73!�"J��"	��<�j�M
p=;3 ��[A��ݨ�S�"I�TN%���I'9�S4D�$������2ky�k���j�ʵqV���ٽA���I$�|�����)�3�m�td��dr�9v��q�����9�vL�18/����I$�Kz{��vU��Vv�\�.�K\���s(����ɻ.:ڪ�K.�I$IYYy��8b�y�8����6Nщ��$Vb�(��x�cJV�n]?�, p$�H$�$�� 8N�$��L(K�FK��V�uc��L`�6`�l`�6�6�L0l������l>p�1�6���,�	h),�	�%
Y#�b��aZ�%�TeZ��7���m$o��]w�:V�b�#I��za��{��_��hz�^���׏;c�R�՛[����x
/�Ϗ�#��UN5~%����E2c @�1�圯*���t������ wChd��J����ǈ���'0��M��x�)�)��ڐ<�f����������^�eobd3r��b�쨭E@�Ѫ�]M�k7xo(m�z����9�s(�[F ��D�� j�I��<�'q1*Q��I&�N,���
�2�%ov���2�lsT.1^��+ִ��.�������� ]r���)�
�;�m�W��c]ڂ�q�Y#A[�?���khF6�w�u�@"n*�(�Wp��<s��:�K�{� ��Hj�iy��P0O���5��!ľ�v��?6U(	 �C����,/��P_��'	��(����[��ʣ���R�%����HE�3�������6Y �+���7�";���@yeTC�eW��9jC�.i3����Yf��7P#%��ںHH ���Z�fV'�f�L���4Q��Xf��A�¹���o:��),
d|�zޕ�z��)y�`�R�Z�� i>S3iH�ۙ��(IKH$�SUœ�q��nJ%���p<��5�y�(N[Js��;!�ӝ�� X��dѡO�T@� �l�h��)�F�?�