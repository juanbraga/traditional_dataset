BZh91AY&SY���@ 
_�Px����߰����P���f4C�Z��m6$�hhLL�mO�&�L�#�d���4�JG�h1 ��  "&���h��)�d4� hhjJ���d�L& ��d`0$��SS�G��Sz�(F����z 2 z���	�y�H���	'H��h;hyՔ0%��s%��{�./I4�ch���5[]�.��p�m��q��HoaI�86Ym��"�Z����3]*�6�JIR�՞u1$L�`g�Y�������92����Cu�W��ydh0���z�o)�����L�BA�m�lc�H%�0�Wy�5�!��^s�Q��2�Ӗ�h������qp���2u� �0͊Ya���wv|xr�P)@H��2�!͐�Q�@�T����	�v fɈ��g��۴ �¢�Yk:��GCM��n�>|�F'Ut��gL�+*���\6�����\���̭k`�\V��s���0̭$at6�˰�����BWom/���B-ڢ�cUO�2�w|�i���$Z�`1�Ů-��w^�I��66���`�"'�˹O8�����*�b�*rV,�g-��\���Q�M�"�h��p{�%�Qy�H���9���0����O�bHŘ����ݔGqDj���k�r]k������}����W�w��x#-���J	u|���g�.���TJ�(��y7t�����H�d�Y��eq��+=�t$v�M��z���=��$����Ci��p���Q��m���Q�'<����v/�u�~���:��K7w8�����e"���E��#Jae�J���=�I	��B�'���bh޼�\��r����K��+]��K�i9P�k|��8��,�Qq���Tj�\�8�ϕ2����Aj�#�ۣ�c�+��M��
,l'�W�D@�O��$�G4�"jjfS���)�Fq�Gl2��X��?K#�R8��*p��a�Locbv@}kDr�_>�ZB+��2a�����mӎ���1�R��i� I��q�Za�m��\L0��,CA�(�	ɶ1����M�$(�U鮒PrJ�y�' �l"5�F"�UY�U����L�ԍ���2�N�v$=8QrB3�'Aɶ�䡶ߜ<}��4�.�=��G]�aҮb8�F'9��*�Ɛ��n �p,L�Hf	��;$k)�%�W_;VT�l���e����R���^s����Xq����� �dȤ���5ju�5�'1*�d�@�lSc��XÂ+"��Ql���)I��>��-�*I��"'<L�V��!\/_�g�g;ՇC\�y�6d����kSE�>�xq�1��<C2a��pU�rE8P����@