BZh91AY&SY�)� v�_�py���������`K  ƀ(( �    ��;�6bH��KKj"Z�J � �`Th ֥*��A+l�Je�R��"�-�Q6J��E-4�Ib�[d���fEK&T� �T��B�#R��lT3j���    j��@J�2d�45 �   "��	J�F  !�&�  ��db0�`!�M0�!�F��j~�T�U)��h�2M2i��@ i&��=C�h @ ��  D�@��i��a�b�����MO�S�����Z��,>�UE�n��)B�+�O�U���?x~�~��FA���Ơ|��az���uE�� h��{�TA\D�>�GD�=?W_�.���@	$@�BE{ �F@	 d�H!PBDI$I**TVEd�B��� ��	� ZH� ��x%ॠ%D�%Ad�D		$T�D$D�B�%@d�B�Z����P��"$�,�ȃ # ��%� Z"H��Z(ZH) �"Z"H�@����TU� +x��U��[5Ԧ�Q�����p�M�Bե��\��w�l�ZLi�B��jZpe�߯[mI�j���v�A9xk2ST�Kv�i�k%%�4T��'�g�o�SQ+���Y�V_]@��Nȫ���#�d��a���MY���M�-�/#��`�b��#	f�]!)�e\6)�[Tu,*�e��H���X[j�Ǹ	H9YZ�ni�!'�y[�fhR�y���f���V�-n�\"�1	��am#cb�I��5��/H��c7j�V�����=���cj�ͫ��*e�ٛ�]�H�F��U{���ٺ���j ��d�S�;�G�ێ���;F�V=)&�:��S�o�p�j���x$�)qJ�o)L��jL�L�NVc�ب1�� ��Y)S8���n)v+7e�ۦ�ޫ³M<�HJ��{Y{`ař��Pմ�M�k%Ën#��`X�ri�f^�n�h340��/Sy�M&/�'*�KZ	�`��a�G�7���Z�;O.���l}�[��!j�K�kw��R�Tr��<NkTD��2
h���3�j�=�j�hkrQ�̺�)8v�Ѡ)m�2=�˹��8�,�w.�N��2��ٲ*V)��M�V͎�l��&��{�Ye���3��a Mv&�D̷w��RE=N��Tn3h33r��-���W��4Br-zc�R����+x��k�95a�ެȖ��[���kmLO�[/�7u1f�Yf�-a���q�o(D��u3b�l��\�������F�8z�|0դolf�%�"�A{)C��C��XvMcu*����Y���0˘H�F+Bt�m���9�X+&���u&�U8TE
�V�	?"#Z����WmhN���:3y0o����-���[���7�}�����Cv���%|�E��\���'�}?Lע�<r�	M[q��knn�.Մy���M���M�VY���)♱�-��v�VYHZ�aa5f����^kt&ц�+�V�k1�-]j���7����Z[MGr)��Ru�u�M��lY�9�k��mBŋ*b[sÚ����2�����UHa����cl���h���3A�u�0հ��[��t���n�8lmu��旅�)
4Κm�]�t�n�+2���n����,q�M��.�F�f�q)T�39��V�%M������w5��M�ye-�6�Yj2ᤪQ��(�
٦�j�u�:��[ "�VT	uW"qau[Ths�-[��Y��J4�B�, �Y����:"����%�Abk���iB�ƕ��� �ݒ�р\9&�kY����l�������2�m%�Y��"�`�ҲR���K.k��9j����,��kt*KY�)�V�[-5k,3	n��r��qͥ��Y�kMd��e�j@��]=G�n��]m+���ձ��Q�M˴-�5eĥ�hh��jKJ��s2�V�-�´#.� *�n�e�bE�-6�+��o�י�X��X[��mV,ܴ��]5ef�.[�ҚP��s.�2[˶ԑn�a��Gh����J��\���\�u���PAy���ࢢ猷\Aϋ��Q,��N\շ T��G�]X(����_��ר:g�?땸��"y�gVU?�������R�3��ص�m!��)^���\���V41��H�4	�z�J�G<6ʑ �)6!0b��5�l����bf�]lk�4��81 ��)���n�.��a΍ֺ��59�� fiEMa�Rk��3Ź�Yc�Xʱ�a�m�,�6F[)�m巚;E��Ԝ�$��9������~�鎋�+f���k*�ffܕ������\s�'�K���M�]�mkV���JL��LSR������eU�k�t��dRRIUEԭ��h�c<���(J���25��V��קX�jP�Y�.�겋Y�{���D/T�����kd��-�g2����*�2�i1Kh��Sm��|�<r������zs�tNN�I H�g&9�y<�u���w�+�]w(a���D�O�F� �)���u���P�dDĴ	$�X� Zc:_k./Nz�Ē���P�j�mE2B�k�ؾP�TFMb�*t��i��B�ɡ%��B�v�ɵ�OS5MԐ$g/�τ���' ':#�~d H˳I ��� Y5Q��$�L��r�#�������\#{��c싺&��#�>g�d�?AUy2;(�#��@@� s�M��~���F��q����8��a޹);%=Ò �Y��xF6��}w��;����%��5%��/���ߗ�D�ΰĄ(@>���^�/��T&S+&q1#�H�Ix�A#���5�N�D�v���w|���0���\�:`��	I�+Yjkn=�>op���Np<�ê� '���sՔ H��|(R>=w��;$�OM�ظ�i)��{Z��#�]2$���Q��$dI�0�
�����F���8R��6ڡ�Y6��e�dK��]��V�0���^kl���g�9�I��x�|ۗ'��6e	&�B�. Ʉz�������܁D����V�b#H�������	�� y`�Io!�.n�ϝr��������]SV�����1�ȒiTYɯ���&H�PAO"�T:�'�t���D���؍���&.$*&]����'~ �"���"cwo\��4&��
w�V��r�&�!�7�?���`���J�ulg�+�/�k��>E������]����s"����]*��v���=��c"@�7׭պ�h�w٩���ΐ�EAA�=` #�'�j~eJsզ�͎�#�Э���ްJ���c5`����G�{;>�::-��
�d�PJ&��1=�$���'�0�C�[��V���fPh1�Y����P�6��3]�}���=��u˺�#b���f�+n���ȀbTI4��c�VT͉5�+�V`��a�c�9�g��oO=���y6V`�n`�tb"L�#2Wg)&�.~]��;�_{��c�v���~��.I�.���V~�H��FB�����#������1��s'�ge�����5��y�,|��F0�y����У'��/�(��Y��2t��
P��(���q�(��ST"!����}nNW?����~2:��a������U�� ��N�rs�B�f�Jඖʙ֞a��l�+�V�!3�ggϒ/��H��h=�����ÚK[sZ�<>��D@�a�o��?@�B��9����TwL�8���+1��B�u^����p���U!D"�Q�ʷ�7I��YN�x	��K��}>�<�"���6��a2����89��TfބM-ML���!�zc^�?-��)��I�� x��\3l	���Ȭ�^��J�PY4���x��<��1��)/</h�u��(==L7��{w+.r$����{����'/��4���&��%��K�F�hm-H�q����p������r(�XA�}W�*���aH#�x½����T՞f�7*�ID4�e�öjEu�١�?���|c�6g�B&�s���^�7�!�����[$f�P�� �O�њ7U��շ��ڽ���@0a�B�'�T"`m����35�|�D�N"ǳEר0tu����~_���?`���۟��2�~[z<�+}j�nTw�6\;ݹ>�g��s���^�ѕ�{�鋊J1��E@��!q-�f�?]�y�1=�e��g�<�F�� ;���~$ \���)���rJ^�)O��s�k�%l}�;"Z����<2oǺ`�,6��'��F*���[>�렘���G;J'�"����P��Əj���ʜ��g�%�]0�@���|��E`d����:>P�2�b�f�Vh�0,l��9��e}h��~�wנ>�Y�a���tde\��"z����Z��]-/%eu1�^?c��c��ꭑ>����0=��"E�?U{ӴUEq&�[�⚍��h��dH�G�$��"Λ#�?��M9����]N6&%x����Xi��5�Ő�@jF<Y5����J���^w\����3%zM/��*^�\YN����?l3�)�(�s���A*����w�<�A���f����b8��GX��=�/=g����!ݳ�<i�T��|n�0��χG��p0�f����-���'8|h��`�չ���^��z=#0�y�u�nCp��'�y�("��V���{P��e�#J%���353��Q}0B/FJ��L�D��CL%��z"����٢�L)'tk8���#dd�ȝ����te]��}t�e���{j=��B}���*r4g��4�6!�	+���02Ю�*�����
;R�F��WV��T�fs�X�K�����i��M�F�WDLٴs���t�R�f��9`��Keyr�؎tYh�Jݣ�aB)!5��,��lP�>�G��W�w�{ăD���LH]u���ɶ�#S4v��e��h�1	�b�������Sv*�~^>�ۖ�5��wU�??T���\�鱵UMH��s�r=�͑dcڞܓZ% oS�ǫ�v��ȧ�ժK+M���`�=�e�k(Ux�9=��}1�*�p)�
����TF�1�h��I��P�0��K+�;���z���¥���Df�!$vݹ�Z�r��9Y�o�p����@���J�k���À�e\��:ja!7
�&H����]���׽Y|*;&gƹ������!N��j��^��/�G	�v#ju�$��6h�)J�{�B����'.�����tI��Қuc���_�ț�]��J�ULx�L��}�j�Z5��s.���N�� D��@�=m/
B����Z��̀Fn2���M��M����z��:��0렷ޥ[\��^F�l��o������a��j�굺�P7�RQ��F�[����D�:�h���e�����[ڞ���p#��,�[O<�x�E�����c���)�q��Sm-ɽ����ƕ��i�A���~+c�����?G]�r�׫�~ �^��n���v��XbM;�LDG�=�3�*��#2���l����O�@�y�=�;dz?O\�������=�O6�c�{�k��3��U�_D��4�{��L�i���~N���H�,�"���d�*h	X����)~�
z�Z\����;�E���֌�w>�.g?�Kƨ<��徊��n1x`��'�B�%��M6�LU�E�f+�ܣtf�Q�yv6�ƴX��#qh5<!�C��}
9����p"2����9$���*��DA�YK(u�]ND$� [���%bA���C,�����3}��&v�C"����yQ>�=6������g'w:�_o�lC�i;���a�7ˋv��n�/�
M�L"F�GoMtZt��g���Z
�[�=��\�sS�{�<�9Ο�a����V�|i��)�cv��U��7���GBL���zwf�jp\oz����&���Z.�%N� �>�U�\�N�7tq�}�SJ�2�X�R�J�z��M�Ǖ:]��R�i\o��jaq�:cO���½}̊����-�����,~1��i.��r7�^ _LD��?t��u�'yj��z=���v���<�=ѕ��\�A %, �$��Fy��,̰���-��3]�#Ư _��i¥�֢n�����t�y� �Fe��?D^���˞��4��0HC��Է��K�Q����'k6>�+��ʃ{�d�ta��
Ԥ��t<:H'��6�X�Q0"��	j	ZD[�;�~��ݑ>S�9uf~���T=��u�7�� PHN�W*�v�i{i��M=�G�5lv8�P�Qu�Ճ�D�s��*�]�Q�'g�Nz��M��6�Юq��5��|��c��ug�Z��m�P�unT�Y�V��c3�2}V}:�_��#-;1�ِM4#�9����t����Q��Qa�%%sWn«z�7�;L�h��(*W��9�#�g�&V�h;�i,�^�af��3�W#����)���uڴ�%qjo��V+(M�֭��%��.#�]�k�Hk�{{"qu�J�v�P�1��,���!V��z���������7!�����W:�8Hk

0_W}<)�|��_1�����k�>��sMlG����pp<�s����D��;��	][mqs��*���FI�����*s�JO(`"z �j�qx�tj�`��Ӹ��epkĆ.�q��bzɁyfo�x�vb�m�[�	E ���>�4M��F��˒"���Kwu�4�5ҭъ���r�!ϐ��~���x��$�����g������:_�k-��ʫ3.ڏ�H�%Ҥ��:\̄�G"$����4�Z�����wh�ewס^ҹC::Ծ�piu���0>��r�h���8�Z�ɉf��F�Vе��l��m��B�[��R�@�j�0	Ij͂�"ۈ��j���+��
B׊�sp��ʄ��Ԍ���c�-�xB��CA�rR�)�r�Ԇl]૴u�r3�/��:�������\�Z93)pg[n����ж�nx=zyĶ1´�r���<�+��p��d���'2��˟f�����ב��z��O yD��XIPK��Ļ�΅��?)��D1�/p7!{���=N�K�6���wuS��SP�!�ѥ����Eo9�����
-���Y��b]"�0�-3پ�ho��s]��VL�td���۶.����7�}wZ'C�����'2�zk��I,=�b��~�m�{�	�>��p��ݕ�1W!�0K�6�x��뉦� R��m�T��k��Mߗ���C�T�;�]�U9�<WF?<	^6l*&��fN	�k���̌[V4"g,��*lS+r�n],"͖�V��H �V����U��DN����\�Td򲨹p�#yN�̳8Q��������Oլԉ@*JT�fR���7^����o��2�S��ɩ|��<ۧP��%�/_��귭l�nP�c��a�6]C�3�`���7���sne�[�ξ��+%�=iumA\v�A��mTt60�D��	�;�0�0-���5��)�<��8;����~ᐟ`k:��{�?N��h�U�u�|���品�5w�mڢM"����a%\��/�P�D�罻-��Mn��'iEl[��9s�hk�C1����ZS���n��(��k���֚� ;�Ң���
��_6���u+yח�����^�MѴ]�|ˣ}ʤr�v�ۛ���,��Y0#�K��u�P&#�v��[*��ZH&���M��v�JXB�0�.-����a%eQ�3I�#����4a����8\���]ɕ��?������/��4 ǳP����E�1K�v.�����_��?���Y�Ն	��9T̸��J"b�8�ō�e�ݟ�RV���p(������ڂ��C�v/�	�J ���Ay���8����B��Ff��)x#��ׁ�?ͷ�<,��5��%��{��(u���{�S<���S�����Տ��Gra��r�����R�ޫ����%5�5F me?i"��t� 7�L�W��P�/w�n��gp׀����>��3}ŷ[����$|>Ź��͑�a��Vh|>m
P�0D.��k�r�l�%A�5�vR{����	�<B�ꕹs"��x��ߜ׎���槊T{F/��=���iB�]W�h�|�y�-��^u�gxlv_Y{�c^h�����g.�L����ɜ,�	�K%%���ˉiqQ���SN�h�%mTdOK��Ư^>��'����e@�+u��X�44��  ��x9�o�\�n6�����K~��ZH��zy�=�Am�S��r^��dzπ���>�8i��"z�]�J����GVߺ	�1VyC��",�l�qx�n���1���p96n�;��"k}a/�I��C@.���;[�f�B;F����5wU7��-Z�5w$��8��� ��]���3��f�(���*�z!����5^�1Ē�ҫ��bg��^:�*;�ZW*[Ǆp(�f�ላ7�:�
>���&�r�h�F ��l���tH�:W�'���P��Ck����/h��f:f8\Y��Gi���r8�H��= Ln���C4]֒J�T7�$�Qq���Κ!Lgr�X�{;-����w����6���v�3{M�j��x<��j0��h��1p3:�t���C��L�����:B�ᰮ��7!X۹v�MGO��~���	���7���G��yB7+b�/He]����x�M�rny�1뻾2s�f=N��C�r��wJ��>[I�Ѵ�3�8��}[Yg��Ci�RG�7��(G��Y �a�ًs�u�)q�5�l��e��]�ږ�	��0��ű��:Ԗ.��,�x��t�q*�i�5�k��m7(E�Ա�6����V��d�Ȑ�NPr�G;]�K.�,�Ɗ-����q�S\��r�_GR���[)p�"�g��^hd��$�al3ۺ���MIF���kE��o��Ż�nm�Q@��Б^+5/s�y��7|6��;���ƃa����������Q�a�4���n����o���^Wa����"*zw�������i��9�8H���hzh�z��1)O��6I�=��ݎX�
��sk��(�r�n��ǹ�F���+��h����Y�3=����(��F�_A�ڷ�)�N{�G>kj����2�֎ܳ*����G��8&Ґ1��{u�u�2g"��m��՛[7}��3&s�fh��&P#>�Ⴓ�R��@�! 	vB˴��f���ʏ����.CA���L�����T�#���̞������2�,��"	mh���`�{v�p�6(����� �M��`*D�Tpy������{bl,�42P�*���S��h�Wou�.S�ʂ"tJv��;׊w'��������y�ne�{�;�r�Gc�E��ko�>�k��j7\��G�e$�f#nml�3E��g�{�xH���>��`+.���^�o4-���e�����=狎	^�H�%YC7Gʭ�ўЯ|���Nv��X�O۫���E`���:|_�*���{H�砧3�
���R��6�ats�U��f�풃tl�DU�*��^�T_i`��y��OOc:m@3G��{+ꉃ���+��R��l�/6}T]f�n!��*6L��֊�޾��GV������l,�N�E���*�9´ɨ�ɭ����R�m�p\���1u|��#�.���B:f�tF�"�9��?��ʢ������W���G�-��,ƤLv��;S�E�v�{��N���+ge]��ɸŭ��|�#��slN�Gm\r��4��)���k�물u�����Y�ų廐^O`�̂���2����D�c�Ba�[�y�}�#��T�ϰd7^��:��ܲ?�:��O�����[��=*n8%^�<O��e���;��_���®+1yR@�-"f�0��?!	�t$k���6���}�z�w߳׳� �n��4ym����Q�"Kf~h�SU˭Bw��  �|�{_����گ�k�`.֟����pZ������N����&���0��^Ovb˕����ZT�N2 S�nED����F;/i��P�!��������΀UeU�J�:�2���dz3�4�Q���Yx(^�ebA��}�V�[�s|�A��K�j���8M2�n��#::�p��)vlL���ޅ� �+��㊼�`���9i)���9�q.�*b(;�Ap�
�si�:���.b�i��zT*Tnꔟ��ٍeߢ�^^��w��y�I�YYSgk3Eڦ�v��Q�V̺�L�˻��׽�x0^iV�7��cj��������>)'��흯�M�}�\NwU�����\L<Y�a�g���%���9O��;4�r64]u�D��l����
wg���4�ͽ��A�Zh�t�8����r'6�3%vU�����T̽"�%Nr�����A�"�
��ȷ˪yn1d~q{]����^�Һ��i��T6���5N{��������Э��� ��eګ%g�/w/D���Ki>
���d���Mv2Ǣ���N���>V/{!��cE��u��7)��ԯn�����^�B�j��RN��,���6�	�~{��TN�],;v����7�AwA�v��g�l���f���3��κˑ^��(�h0e�3THn������3h����[x��%�n&���Rg���x���7��+m1��mF�4�,��4��5�!l��s\�Dˊ�n[�pme\b����X�ن�f�:�mx�Cq�5Ycs��V�+5��ԭt�o_d�\}�h���f�	6�X������ᔑpS,��[�İ�Qm�E�]���m�l�r0)����٣�� ljq�ގ�$��1p���N�WJ횴�)���̵T�q��\u���Z���z3�]L[�Lsn'���Ϗl2AإI|P���7�D�Q�yԽ��)�p�kz
F�}�0���;�m���Р��D'�Y�u��/mϧx,-��y`${u�s�������nd-]�x��7Y��q]C[sgX��6�%��4��q�ƙ�7���뿣�4��}r���>��{՛O�hؾ;*
�6�蹶�%��S��n�1�[6��(�Җ��HI���y@�j�KpS}��[�;�L �Y��Ҹ�hwq����i�2��d��u�Gԍj*v/Zx�[㉾��#��y�پqA!��"�o���sL�J2���v��=�i�g�Ǻo:vu� �����'�_{l���l߼����h��~r�v9R��O���k۾���:�J��7gΔXXË��QU�fC��.ŷ�w*"!\��
�[�s�tr��>9��@�X����@��w=Ҷ-bP�ج��h�;=���HH�����^ RuW�4�����p�uJ\�
kw-�Ω��m*�B�u.:޼���tן<�;h-��y}�c6i���Ku�Rj�8F{��ސ�%��M(o�.�s���Y�ﲒ�h�Pt�uw�m�be\X53O�����K��V8��㝘�u��sfx�,�m �׫5/n���=oz�Z��!ܮh�����9T]�'_f^ZRp�P��7�e)e���ðWy��L���%��6<��vQ�$Hf�V� U@���%h\�b���%����.����몀��+����H��KP���܀�u�B�7r��#�4ڄ��vY؇ƫe�S#*�^��1���C�FJ�v�nͮ�==�i<������;�9��AR���s7���)�+�Kz!�y�@�^�J֎�з����%��g���]6��Yq�KX�	�S2�%̣a�H�%�0�ot���:>yM��Dp�<����X�|�1Y��-��oy]:�L-
ET�s�P���0��*~�h�ݻ*,��������0tlWd����j+"!P��ny�l��L��w�'��Ҧ�I��k����Ϝ�9�<[8�%d&$[ہ,��-�`ܹ�/y*ʤ��g<v��t�I��������heB�z^g[9��eԿ@'u�m�.�@��u��k�{�jO9�R�=�">��|�8e_
�yYT���M[��=��_^�(u��Kct�&�R���m�\SVn9����d檵<8C�vh�q�W�/t��>����w���N�x	"�%�;��2��I�:�1S�',�7������������6�M�Z�ݳ�v箵�;�1�bw͸D���-ln,�;9��S�$cdf�� m��+w����M��s;0o����ʃ&�T�D�C���ndI�[=�О1�/�zfn��gC�Z�T�A��Q@�!��^��?NA��k�Bwk��^ά�P�%gM��t�{S��~_��?����H òI"EEE������{Og�/��Ƿ��a�\{�rD�-��!h^��RDE~PA�ئY ��AȈک?�*-(E����-�
�EUA �$���*^�|�e"k^��|(7A�ΓX�����$T@n��H�cKL�e)�` ��Q�-0D�Tt��E�u0#�A�b����M�]KnԖu�'����zӷ>T�V�u��S��}�K��o%��6�W���u�r>`QD�<;����ۤ����zο�����ĄT_�*I)����=�ǟ���/V����e-���~/��!~;�r��y�?EE���?��]�i`�F��`�����[6��D�T9�X��\��i�f�N��9{!醙_���(g>e���.L�,)-;��-� �
��T
�ޅ%���Q�w_b�]�f������ȁNQ
Im�n|�X�9�ez�Bk�tV�B���=፱�E�?m�����B���������c�ʊ��d�r�g��m��i�ӧ�ȟ_Y�n�=|j�uw�F�z=���������帼��~��Z�����TdbN���'��$��-o����mv�a�0��y<�Plw�*/�}��NzN�}Y��O
�Y,]6'ī��L���B���\�B3Ļ�Fir�Pi}r��#�.M���bQ6i�?�IOnB�]S7���7�B��lZL3��
��d0����j�����N�EE����9�e�L��q7�0����׀~:��,.��U<����H���������;8�Ѽ ���Wf�:��BҐ�o�s��EE����Vg��i��n��>�r���D��̐�]�N�&�	D���p�q�nhk�:�۞��\���u8exe�.�o᳑͘�|�QQn���ۦB.G%�[�)�f���sp߱�x�o�Ne[�������x9���8��E�/��C�^D�Cu����ft��P�s�J�����e�gI���z�'�z:-!�U#�c������]��BC�̧�