BZh91AY&SY��Wq �߀Py����߰����`?�w�޸۸��$Pp�  HJ#Hz)��ԟ��L�z��OH�&����@5Oi�Ҥ� d4 ���  j��Ri�T4  22h � 5=R~��A�      �&L��L �0L�0�RD!�*~���4�'�L&��1597bH�2Q%�BZ4���/KO����^��D��j���0��Oفl����J��(B�B���6j�|v<�#C-�6C
iB�!1�h#c�1�hl�cA�hq�� ��T:�=�B�e���,��,��,@�Ym�YIB�kv�ke�Ye�:�&6*����F�V��r�~�l]�@��m�2��%d)S3"��U�R�i)�>���٫&�;;*	v*1��wL�U���e͋Ȝ����a�j0�;qA�$c5:,8(�k"���vr�w4�r��ip�v����gv�q�����lm��%�ƜQ��G�Ҩ����]�\aGbRP���tS1�)-��Za���me���Q8��:b�+��	M��)��x�䥫;��/�]���vvv��gggggf�i�:�[oi��r�Mbi��M4�M4�o[�m����Mbi��r�:i�������r�:��M4�N��q���|�u$TT�[��szN�MF�G11��
��������Te�F��qj����E`B
���
'��U��m�_�h�蝟�W�H/V
:"a�x{&:Q��b���g^����&��
��(`/#1D��k� x ϑ�n�����X�c�����    �T�o6�u�Y�C�g9���"j�\W��yG�.*�
� 8���c4�<��
�"H���{7 Yy�6[>	������f׭��ALnG��o:��\b�    p�>������RSA�YTr6\��8Rј�@�pu�5P��;�$�ܐ��q�����(o�@�غŗb6��R��q!*N֓S���
�c�K;W�X�   �m6�=T�u�c,w�̏5_]D�����bs*%1;�Av:r��E��v(t���b���2�n�N1�,�9ƚU��Ur�:�%����:��g������sw�   <�`�	Y�����$�����S�=�6c�=$@D iU&R^�{E^��w���
y�@M����*A�KD.}�6.����I$�In$��qݙ1�Ҋ�+�@R�Eya��=��}���켨ˢd�q{S�b�=N��:�|EUL9�q��^q4�{�f2j�(���,�   I$��Cc�O59t֔bNG��E���_�C7U�]��\f=F
��D�&@����35�r��}A�sr|kz��˼i��ֹ�   y��Yr��O`�2�toU��.Xjn� �9��0��tǏ�ś��ȑYuBz-�$J�9���)��y�:~Lf�@  �:�y�|g���{�ۻE5��i�垑�%}OY<��>��IB̥�J0����ٳ�TR��Nރc���1�S:c�V�\�TK�mJI)I$�f^��X7mC����a����G�ɑ��0U��mM\4®��:��7�}S���-*X��r�
[�q|	�x)JU)U�UR�� U����������&O�n���R������,QE(�¬T��)ER�U��)��J(����QE(���)EJ*QJ)ER��*U�QR��R�c䴖(��R�QW���/K^��\JT�,,^䗪��֘ P�ь��bسU&*2���9� �I�뎽�j����CZ�r�T��bg>(i$j?7�4/ۺ�O��6��Ɠ6Ǝ�ovθ����]��mw7�e eyg�r��^Y�ϊ�3]Wi������%M��H�?����y�yh�7�/���ɓTR��ZR����H�q�^�l�=n��1���d�ZLq��b��=	Ԑҩ�;:��g'^k�žy{���)eG2����Oe�{��J�j�-��{�ύ�i���wᅘ/V�7���{}�`BtJ�!��ii��ͺ,{4�`�dx1��?�"҄������k4�r�I���u�������,�NI��}'VRb���l}:i��~��:]=>*X����c��s�-.�ߗ\~�G/a��ɡgE�te$��86�Xγ�q,�-+g<��#'t�F�ʥQEr5r,ú|y�K-�8�g�M���"����=�r�u>i�L$�)�)��JZR.��cF��6�4YN9}�3H8��w�1��i#��%����.�b�*~��&Q�)�ʪ�Y/0���XL�z�4=�R Z�)1�5q�}�O�%vs39�$J/#���"ﱆ��{$�y��{��H�5���*��oQ)�wϙ��R3�*p�@Y��`EԴw:' �Y$��$��^=>�l�}��&�=�[lo�K8ټb�ʲl��;n阰�|"��s��_~���M��{g��I�g&�f�s's��C4�)���� 1T���9&��V����[{���^(�D�T�*Bگ��(e���1)2٢A�P��[��n�QH�i���M\����:��;��*��:f9�Y:*�zeE	�K�]?���)����