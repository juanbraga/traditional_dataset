BZh91AY&SYb��
 =߀px����߰����P�J��$ �"hM�F��L��I�  2d�j�O���h��F� �����I�Q���#Ȧ��ѧ��4ɠ��zC��2b10d�2 h�00dɓ��&	�F�!���s%f$JJR I�z�������̆����D���ml����b�o)�����\�c�}�J��Z�ʑ�ӰƸ��Gp�Y�VIS,ǟs�{�#��2}&['�b�Ԑ��) ��u�^���M7�xw�y��f_�.�|��[�+<Eas��dg��3�? ^D�c��Ug�PR,`��Z�QPp� ƥ�ٕA��ţ������llm�6�8=xs)��]�hQ�U��x����1�>9�?�R�3�K�����
��U�-�R0�$��
�V`f��ң�ٍ�ӈ������8>��ޭd��5��h�-E��r��.�9�:��Gƃ�~T���n��g��Q�J��fI׆�N_9�?1��E(v'����"�#����3	x���B�����!ep#�8N�d쬒�afv��
��d��_ϗwV�׊2*��Ǳ���� ��i�e%��ב�h�\�S�#%�*S�zҸ�K�״�8՗��F�A2��Ivd1<q�84b�i��Y���+�Ƽ�vP���)Qa�!g���f�F�#��[��m��X��lc�s�<9UG~���N�p����u΁T��Ri�Q
S\�q\��
*rК������P%&Ȓ�	�g��Tb�*a ɢ�x2���:�:��h�ɦ����B��_9�N��˦�/���8���Ӗ���ʡ��9��<��X��{x�u&Q�gN����ʥ�kgϺV����h�������)P�h��}����.u�3�a��P2�bh^�����CSf��3l�(�m6�F�.ͅ���,�]�򼑮&a�(6���T��+\�*�QJ�dt`3duۚ�e�-SOl�U��L��x<���rE8P�b��
