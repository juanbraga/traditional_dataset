BZh91AY&SY�I5� ߀Px����߰����P9n�B�'Z�	$&M4h����mA�=&�@��A�x�M    4  S$D��OQ�&�h���`LM&L�LM2100	i�2�7�Oh��!�� �2	+�	
��I �	�܀_ߍIbGj3]}�������m̣��������͓*q��C;"5�~�x��"w�p(�8�7�6T"U	t�4i�in��͜��hP�M���8��g�L�����E4�@'ee �����Ņ���͗4li��zLW�v1�q�h_mb��j�����J*M,:Bn4�,F�ae�u�v�1h1g3
r�\D �QG�!dɶ'������ή�qr!AE*�t\EV`P��5��B)L�����qRM �Yk�����+��bIzK(�����plF�NB��IU ���)t�"Z�D*dҬ@s��	�NW^��)Tx�gyz%}�u���3�^l�޳�����RBBK�$���O�i<3C��0-�����H�E�4��@_��5a@]��2�It�!G�Ea5\لUE�Wê�
 #Tm��<g���K�o�dt�����ݗ��w���uZtu��Ʈ"H�ɭ���٘@�n����<m%4������3���&��M�L�\���'��2�$6�]�fC�ua��l�/Ȋ��7��(qE�/�Aw� �cm��X�jp�r��j)��.����w���N	�J6?)^Y���Eؾ������H�Я%1�,�!S���.F���Z8�h
�9H2t�gWg�����E�r�@,e|�+�
�k��2% ��X�fs=lC��u�Ơ_�v�]��v�
���]�P`Z�	�Um��cix�Ye�̘gO(�l<s�Z߈�)�`BW�G�s�]���,�\�U�Cī(��(��5$BL2�9�MK��R!�č��{�>�b5
�:��G%@M�-Xn*"��X��~�>���4R�\H��1jOꅅ["�)�7즓)!��v���Y�L�m9�R�Y� w�F�1/Y���Ͷ18WH��^���呑fb4=S��Q�)u2��%��F7m�,�Q@�T��A��'$$j�$��N(C R��|FD�8*b�J�i�̺tΪ�?5uԇ���x�"Ր�c���%r�\�Zj��&���u��%+]6d�Y2Z�+|n��.�p�!��kf