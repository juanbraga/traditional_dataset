BZh91AY&SY�g� q߀Px����߰����`~}��� �>�U>�Fh8I!4)��2ԏSC���ѓ �? 
�C&L�2d� #C�0jx�4�C!�   4����@��1i�4i�� H�H�4�i��   �	iLSi���S�h   4��Q��
LD@�id,|�ڈ��P�p!�D`�8�z�O�@�\i+1�s��Xf/��p��g�!l��A�S$���f���cll:`��D�����d6�i0��110�B@��-�yU[�  �-���u�2�/�{�#l܍FYn>�3!�Ir���G��������$!3&Lιr�;%�����.����n�y̡v��/�����
��IV
� D�=�KʔTJ��%��.� 8�)�:{YX��H'��Z����ۆQ�:Ă6�DV0��6\5%SF�iᱵ�3��ۨi�˘��T�lm�%�
C5�d]��.1�N�tD�QX���[mQ���V��4����X���)�*B�q�����?�ً^�ˈֆ��1l��:q�Rǧ���2P�cH�^/��-�`���I^�p�5b���2�WU�֪۱�ٞЃ%`%	�'rk,l��Z�A�F/r�T�4�u+��^����݋�W+僗�͘lz<��F,6�a�0�X��4��t�J�)��e��8a׏ˣ���q6��޶6@����A��7҂ڰ6�dPX�i'00�K��,J�l$�hnF�Y!	���Aí��U�5^�O$ B&=Ht<N�vv��
]�.���&=nF������	��x��u7���ÿ�My�!E�;�͏�q�j#����*��x$.�y�����rE��#�9��!��/����,�'.j6��dQ+�'=>��!v��1�JB��c��G#��eax:nY��ֶn��7����Jd�E��4v���S�{���xq��LA$�`�Jc�T�K����.�B�_d�',�X+�A��Vc�ѽ���e�t���V�7��A�"�����F�d�P����h��F�j�����V%E�0Z:	�F����+�ݪ��B���cՓ���YR#�kK��re��n��ɶ�[֌gA�ƅ����*gU]AT@�������%uj1K��PV�D�&{+*{60�P�Y��IM�%��$(E�v|95�l4�[�,���fs2O^�VKt���7s'
�w��3�g`�ds[[
�1��#+�jSY�q&�q��Q40�2���a�0��b8hR�0ʔ9�f�Bd8g�=�:��?=8(�Z���u�����*�Md��h�'O����!
������XX�8$�e
VF�V{�U@~z�Y$8YL"�e����]#n���Z�V��-q� ��o×�֧��UF�{&r?�_��H�
 6�� 