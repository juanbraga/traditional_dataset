BZh91AY&SY�B8 v�߀px����߰����`J� j P  =�    ��0�֔�6bN� YaT*$��
Y*
!�XҨ-i �#T3h�L�%$`��+L�%���6b��օIC Z%J�
ٔ%Kl	U�R�� �@��P���6�Tfª�    S��U   �   E?	�)U@       0`��`ѐ��&��OF�Hʨ      F 0`��`ѐ��&��$��&�'��4�LF@4�5=M����U������A[ *
n ����+H������/ �$�
*,
���Ԕ���U	QO�%EA�&��q�'M�B�$� H!"�+��2 H '��B����H,�TT����	 �E	$A�"(Q�BDI$[�/-* * �� HH�"��2!"$�* ���T���EI$ �dD//��E/�B�BAI $@��Ej� dU��@	[ĴR�����Bϼ�`����I�F��$?����>�_� Vd��b�*Ĳlغσ.�ܛ
A��v�l2�w*̕n��̌Y1m]BV�R�%�O)_�jό�T��j��3(+�P���੄n�'R�`V�t�ښ�`-谛���+�b}�kl��
�rYo6��̫)JWz��kx��tUaԍ)\X��	{�&�����V�[�����aA�zFeaSM���Or+{�}��^�1)k.��h�v�W��7e�6%,�ݡ �	��p�Ę7��&Yډa��&���7M�{3t�>H�&�ڝ���9��\
ъ�j��d������r鑑��4]�V�RM�U� ��k�@x,��<�T�{V	W[�8D�2�̲_�RfJ�F�Y����9f�F^'�#����YZ�Si k7`E[�5�O5U�!1�۽��	ŏ32��״ƪ;�J[��ֻ��^�ʹ5C3,ݻt��l�S{���gFi'Y��X�۠�Rp�Xh踆��C3ekim^ F�pس�һ��"�S��&*¬c�.
��,�/ͷH�u;E;i�ܹk^�l�֨d�orR��UZM�[SiQ4�^9/kp	�ø�<���3��n� �E�Nfo�t�/f˭Ю��v.A�p+W,'�֐&$L�bP��J`�3�m;�p�f��%�ͩ�]�dw�M�3[j�w#��,ZnS۹�.��xȉ��,��T�י܄�U�+ۖ�C��ザ���:%`U�)��^���	AS60�_o�Aw��܆P�j�,.^��TCA��J�D*�l�*/�D	V]ԡ�`YJ����(&m�Z�3��z���U��a�;Y�Ro�ބL�ﱾ��Æ�%����v�&���ɉk�ZKi-i$�@�W�m׶==���~l�0��k��X$a�p,ss�՜�7��)�n6v�m��ڰ�``�Sk�3SkU�n�M�)♱�-��v�VYHZ�aa5f����^��M�Ȭn�Z��X�It-��pޭ4�u���wE?�O"yn��D�w6,��5�komBŋ*b[s�kjn���׮\UT�kZ��6����뙠�:�j�]c-�F�YFW7H�lmu���/�(�:i�-v%�m�1Y���t-l1c�Zh5e:�m�m��M�3�[5iBT��ؼ\ Pn�m�k����[��p�U(�cQ�l�J�\��@Ό��U+*���9au[Thv!JZ�9��g@�i�lP���fN�H�1�f����Dq-],J�z�Ҵ���$[�\Z0�$حk6�6p�.e-��⹥L�Ilm�%��+�����F.�˚�uN�H���gW5�%�۩�V�[-5k,3	n��u���6�3Mf��5���٩b�x�5�SMu��@g����j�Bn�B�CV\J^-�IiX���f]պfp�ˢĀ
�[�Yf��`�M�
��d7��٧���X[��mV,�h%6-ںj��N�n�JiB�%̺��o]���u��6�;G�,�.ݥ����z��A�yNy��EE�<��,�@��>�m�o?�Ȩ����EE�HO���m�UI4��P��:�>IYT=���^�u�lR�L��Z+q�S���O�߮�9M�4���SZ�]H獆2�H.�M�L��Mw6W\�S13F��5�`i�����qA�Q�WU0�F�]tu���� fiEMa�Rk��3Ź�Yc�Xʱ�a�m�YJl��S�����-ƞI$�;��~�����_O�c��
٭4t�ʄ�m���%l��n���\?Q�pT�M�@�֭��!m�&�L��X��M�Tb�Rײ��HAI$2�4��[mvѴ1�y��5� m*Z����R�ZR�^�bA�C,gY]#o�u��P�o�$��d��d5�������*�b�v�6�H������*{�:�7����<�3磠t��=��D��&%@	��-F^�km��@V�_	�O�Z�_R,�>�i �$��m��[̶��� �&F$ ���� I�_VL��ޛ�^���<Q}�t�B6���D5�l��i*#&�Y�t��i��
�E�BKb���/�>`���Sy$	���{�_���!�F�	R6�M.Ig���Ah&�,�Gf&!sM���$��U�f�|p�
�x�V�ì{v
p���X�Rͻ�jT���)�a�"�ª���L���
|�h�2�E!��3ϣ�mw���t��J}C�.�M��F6�t�}{ܐ=��$�$�}�q>�_���}��|�M~y�$ 	BI4��^�/K@�LLY3��4���|( ��@�`7���q�v}��������
�_X^^L��^y�������ۏ����<�<���>|<��P|� C�YB��O��#��ߓ��螛	�qxy���qT�ʧ���x��
 Uq��d�i���X�����|@ V��^�^����{��|�}�u���.�i�a�q��^��-qW8Ͽ��X�<�m��>i��C���E���*7GMg���μ���}Fr@�엾��&~i��H�t�����*�*묥c��Ƙ�����h��(@|0|ַM�86��<���U�(E���\�cχ�x=�m�+IӴ���@+R�n�*�i��cT�>���q�����b`D���=i&�B�Y5�tU�^8� �w�*P�g>��}�Ȉ��_��������}�+�_n����YO���������QA8����uQRD�w7:D�L�L����ЪC����´�ӄ�H�`���:'����*۪]�vq@�4��4����ߴW��<�T��r  !���u��L��=ߴPX4,r���2]V�/]c()F�<je���)z�������3���#��d��`@���_۽赸L��;l�,&8
ʙ�&� �aw�G03�t/Ͻ=�w����������b��bs ȶb'D��Xxb�n���X[h ޕL?Z������@P|����D�b�×�&�l�+�iFY�k
����wq1}�V��>���Y��Kޏ��]?Z����f�̵|(-<�b��M�
m�Z�<��SE� C�n��cnYQ5�����1�*��#���a�Q^�UY�����[���~$�ens�[�����i���T���u�����П^V+��fc��9E>�m_r8BG%�һu㧼��q.m�3���￼>�>��1Vw���,TS���Ӡ��1�&g�����FV��U�VI���L2�2��f�A�E){�V�Z�3<>�*�z �������.~lr��0"��iG� ���"3�y�ͳ��eKv��Lk��y�c�ٻV���M���0�4���U\^��{L݋�ܴ�ԥ�X^k�����V�x�;.��7���%G����Wf�e�,(�ۛ��{,r//I̑Ƴ	��)	b�R�Q�	Q)Y �f�4�h��~"�vS���o�E�f�鉲���,oy.6��W��c
n�]X�(�Mp��v��m�q]z�T�琿?ג�a(	\T id�	���7�3���zŤM��/WQ�/�YV�Ӻ�Xz�q�z���� �\3>��FW]Tcn�(2ۯ��&S(��f�z�@��-���ꮢ����'z�9�n���*��\�v��F����*�m���<ɋҽS�{Y���٩��n܉1K�W�l������?��oګp5Sr{�E��b;�����"`'�б+�WL`>��_�3�ҟ'OΓ�Z����O���w���0%$ϼ��D��}y�:�G��TEoK�+�/��V��f QA�l��@���x˴:P��Ҡ�}�Itf� R $O�ȴY�b�f�Vh�0,l��;/�('�i�I��U�M�L*@�%���U�/Lh���=^QsTb��*��u(���4l�ʎ���Z����7���*�7X8}L)���
R�͌���5\=���7[Py�i$F۱X8`�>��JS��de��t���lɼ|;��tӦ��SV�4�WZ�mϸ~�f�L��g�����C��Ø��T�p�֩ؕwK����f8|�iC�)t>~��V��fL�M� m�'y��~M���gFW��O	��냖Gde�vr�ܩ��|��<�L�g06��8�+VcviuvtT�-�cRY��J���K0������^��S{q�L^zn�6�$`y�Lt���9�#�qZ��{�*�7&�fEIk���j�dlwL�\ȉc�٤֠�SN���B�Q�`o,u���V�N���C%�+�����r[3&��`WƘ̈́hr�l��b.�Z�����}��q��� ƙ�f���B��P5�nvv�QڗJ4�eun0�eNL�.bX�)tu0Y���m4�m����6m��Ӻg�m��F�:�
����7b9�e��+v������0"`�B��M�����+~�C>7��]wgjd�m��;J�2�&���ʐ���v㜻�����x����Y���yz�->fBiy�mUR�U"g�?4��hX�#-�ی!$�C]�e��7r9�:o+P���{=�4�P���0�{��<���"]D	�|~z�F�kF��h8�]��G�:t�,�ú�\��b���Qk�2�Fk3Gm�nkfD;��(�E.���ΐ�m ���X�,��t�.�Y�)����P_6�k��J=�׽Y}{~�ϯ=��7�Ľ��)�Nj�ސ�Q�p�I�z��g��b��2����!D�Hm��D	EyG��fҙt��f���w��~�z�>%Wq?�����ݸ?n
O:a4m*�����R�Mn�ֶ�d3s-L&�'I�_f��W*㷶�e���(�� X�n+*�r��E+f:�\��$�I���P�U>�؆z����M4
5��k�r���	��[��\T�tT��̹�;毧��~���s��@ ��R�N3Ԓ��w�{av�
�d'cXC�e>��F��N7�V��I���+WZ2�����Ӹ�j�&Tō5�$�����*���3L�>ܡv߄=�FWs�z�5��0��}]lG��i|�{'����m	Q��
�{��W����m��.���t&�/�ד}ɴ�	�4F�L�J�K`�Z�ȕ�0e�cS<�^��W�������Wo������n��[���4E�#1�ѡ~�o���M���v�mY��7(��e^�]cZ�j5~��*�|�{|}xj5+��2,�ygv�5��g�+!�5���2W��)2��9�v�֪"��/�f�c �=<v �����Q�6��k\��V��X9��FҌнw:��o�bmAPf�W}��06,�ڵ�uN��1R�u(��{o:�s�@�s�ViV��=�.�eW:��p�s��κ���*���A��V�<�b�b��u�$��p��fe	+�CV��V��oPKd���}�R�I9݄�l�ͥ%Fܺ=�[|؉�l����4���G+ J�,S�y���<<���xeH��6B3鼭�æ9���E��oWrO�B���POy֜�^��R����N7�,��/�S |4A֫t���zr��<.G�/:�ɣ�wO�:=��������f�3F����\Us�+�Y�ae��[K�f,�7_��B�@���Չ�����)#���߮5Hw�� x�Z��on5�御��f�%E���m������M}3as�R�8yѳ�s֗+�|�ַ$�����(�8�{�~٥eR\�� .m67��k6����������ɘ=��cN���`�kb�T��!���]�Y����t�.�9?o-�0����(���3��]���[l�hƛ-�A�Mf�WoPє��l_6�h�*L�Ui˔�6�n����V<�x��o��X|�e�l�f�2�b�2�w&��q�9hN��s2�_n��,�M�3��ƊYB��Ez�G;���Ź�叞5sA�}$��|q\�9s1���$����if��N��p�a�s��TՁU�˵��n�iV٪��=��T�޸y"�wTێ݉)r��f2.���f*壞0��������f�p�k+�g��{�#3�J&��ҧ��53˞P�|���D�K���n��>����9I����b	���o����\�XS�Bu�$�ڲ3�J;��I쭡W�D<�a�t|y{�

bVv;��9\(�q�N#_X/�wO)`(苴k{Ŵ�4I=�^+�u�x��	وM�sZ�?z.��i'�b�i�7�Ɏ]0B_���x~��1�n���4}�W�����_eO��-A��Ua�jO�#tUt�}S���!��Ee��������Ho^	��i弥w�KLJ8�����u]e^�dL7��{,n	�Jk(�N9ƪ�vLK5���6궅��#e�mW:jݥ��bU��JKVl�1�F��a����`�!�ySn�Ar�B`�jFk`б�v��<B��CA�rR�)�幩2غ9�Wh���z���ym%�v6�s��h�̥��m�
�f�B۲������,�Fng�U
?|�zg9^YWe�N�.�g��_f�rK6�����|��o),�{�IAKou�[Ϝ�$�W��(�>�tq>�}瞤cȵ xF����]�S��#E
� �D�K�`��ζ���L�QG�hPվZ.n��)�r���o8�:��#��a�1�(��
�{��~�����Cb�����W�-6�w��i��۬�m�==�
��i������-�-����2���9f�j;���nh��W�u�U��M��A��t�˛q�?X%��F霱ƻ$���3nЉ���BېTL�}���c���V�]2���� &h�[IenXm�K�e����m�QN�h�=ICT89HΊ�����(,y`P;e7F�y_Vn�k=���`�ϪF2s�D�J����p�G6C����GLA]��ӎ��fvh�nEK�޸�=~�{of��r�@|Y�F݅EDs9�9e��|1�0O(v���k�[��B�o�ؗ�B�g"+�-��<R�	���8��TJ(����mL{L*�;�n����!o��L���A��u�%�oW6����;Cs�u�����_|f��%M3#Ʊz�m�?Y�`�tq�'���e��0�s����[H�8�{ɧ�s���B'Ӂ�̲|䢎��(��k���֚� ;�*,7A�m�|��J�q�5r����_,�j,�]��Uf��x�eS�C.�{�]yO<A�^e:t��a�X�++h
=�&�!ڣ�Hߝ�dC7Z�`�E7Pn4�4öd�rQd��I�ǵ�d�����sR�5�=~0@U]� b�Ď7l9������>���L_�F�¦��1�+�R��_���������}�z��( �*�h�VET��ܣ���������ؖ%��*L�����w���{:��sA	3WW˂{��<�0��1~=|N�35�R�A�hG�ʗ�_�f��!'�6��ҿ'���F�X<�|���MC�%vmnb�ۦ���Voo"�&�p$j��{��������n�U�R4��N�'}�j����Ĩ��Q����N;3 �y�nz�p�v�n3s��<�������������0d�R�q�!tLkX���fiE�� 2d�`�s]K1.3ŦD��R����g����ͼ����j�R��r��Jy<^�592Q
(#9�y�wN��7<8��t�_���՛'A�j��[�5�wcz{IW�������I����6��G�;.UM)F7�a�$8�SG�|��JK�b�Zpۦ.�p'�PT�8t�M8v�uMև���M�plk��B�V�^�=�=xB>ݔ�R��L�� 8��Dz6�H�E?`x!�EI�V57Q���})k��{Tu�qK3��g�e�3B�N��S7t��-��}�V�h��/�Iҧ�T .�,v�\͈�v�L�<��7륐�2���gS�T��v6�}�r�msu�J��z���$�n�����H]�-�����Պ��Qq�Q��u�$��Dy�JG�}�<��s�P� t�@t��Ϊ��#Jt�vOm
�ś�;]k랣��@n�͞�6(K��7z��H�T��.��;�O8{�� V���TC�I���wfWvs��wO���Hu{j�a�)ea�W�����J.C�ycQU���)g�8������q�|��Sn�*�dLi7��X�~w,��۷�[y��_�>�������}>�\���a"��\g����}�\{Lxw��\����^���t-DU��r�����L?=�li�j�d�U�{/�k�)��eZNI{�x\�̼��y!�� _�i���tn�e.1��������.�mKJ��hbb���jK[�,�x47F�5���V�M���\V��i��^cZ�4�֒�ٙ���qL�9i���Q��b�˄���q��c��4��\lT�#}��=0��V�\�ȻB�l�hd��$�al3��[��&�v�G���<�"z=K"�D&�.8o����U�]�m���fq����-�	B�i�M�%��{G�a�xquW(==��T�vՌ�9[���7�*]��z���Z�SLW2��xjD�|�$�HG�iuђ��U�]aE�c�����Eq�TpW@��r��#7pu���
��rT�^d4�@n���-G3�[scaSyFN}����ś�Ze��9r��y���Z��u{���íD(.�^��WU�vm^�vC�o��b����@L��mi�w�0�y�9xx�5pd��������48��d�R`)Uec66�6Tx��yq�~���p�H�r&a���NS��Ywu��G{VG�X�a�ޓXo&�+3ۣw^����	M�Sj�3�)�}!�=�J�V��mge^R��+mW�:��{ɹ�ta{��j�^�h�7�ZL���eoU��7E��y'xQ�\ԇQ[�8��z�V��|��!�$��$��C\����{/]�T���Q����&���R��م<k�(j���������uЋ��,2���&7�v��7�P�rw5���V�1���t뽨�[H�V�+�É���Ȅ�5s;a�jx�%kt�%B�J�oG=j�"8l�]�[��c���J���ܖgy�z��ii�w&��ܭs�#<O1=��i���|�������t�a�l��듽��|+Ӽ7;hk"D��<�-�NV���?)�3��1F8��n�Y�bЙqii螕%��'&yy�C�sG�Q��5�{���+�8;�P�}<2����y��v{Ye��ң��p����v�\��� ����̲﮲^�4�h�ЧQ�/$�UCwT�ݹ�-�]�����yf]u�buɒՌk�^��	Q�2�	N�S��<oښ��k�r!^ۮ�8�r/u]?�N)Z�p�G=T­x�q���p�^7^�/"Z,����n�=��4#
?:n��®�RGɃ3֪jq���&9u�^튱� �n۔��luT�q5i��(�OU6�m6�fw���Iھ��G��p�b-i�$O���DM�!z���꺅C�dF_;%�� �!c�̜�;Kg藅�b���Q{�wyd����am%��]u:��	0"x��S�'��J�j;qWV+9��xo�i���u,�z��-mNu1�1�x.o�i]�M��	|�)�t���R�w��k�ɓ���l޿z&��&F�F���j98���i�J_I�-F�r��<�,�O+�A��"��O��C�����iN�Z$�B�;�.S���mXK�d`��Or���u�>�n���M#AL�E6��;Mj(�d�fJJ�R�<]��I��(������+)�G�T�+ޘ��I;����Ce�c";����͂��z���9�5r��wxe.�`i����\l]u�-�ֺ4�ig�Y�>f�\ ]L�D��Ѳ.�cG�u����_�������zi�s�W�;$�ɦ��1FeV�����{J�4�.��H�Ϫy�Y�<~�{]��۰��Q��{}5i��B��y��$w�g:Y���c���jC]��*��v��D�2�L�%���*3����OZkm�=J�f8q]B�t�^$����wZ�ŹQ�6P�(��d��f�,��wv��뺒p��φ4����B�׼����FlXs��whhE[�b[[E��[j�Os9�et��t��F6�J(�J�q+� ��$���>M�>�W�b���[y�L�L1����XmI�k��+m�ԗsz��m�3-�Hݵ&���6Ɩf��-�8N�-�2��ո6���1q`
Bܬql�v�MI���Cs�j���vIXЬ��4#R��e��n��\�+�ѵ���,m��MQ���56�L�"�y��`I�������O�ܧ�B[�Mt3Ѩ፦�f�6�=I[򏏈VY@4����]�1;���޹�ݒg��B�ۓ�W_��rm�����:��y�o��z��=�I::o��_ܖCw뤙ME�u�hBb?�Pb��������O-<�-���z�Q������	�f�?h�N�xj�������m�8��z�V��t�{`�ld�/�VB�e��W���)�6�s?�T�[�Y�HGCz/�S�뿇�*o�Vؕ��ѩ�����f���и���2����Ɨ�(��	��l�A0��La�b�KvM��Y��b��B6o*'�n��D����cq'x��+��>ޠ؏���X��I�J�MD\T���&-�B��5Zӝ���3���oN^�:do; _#Q3�&�Aoϳ2��$w=��)��
{uU칲����ތI��v��$����8�C���+gk����E���
��>N��;3�[o���e("n@�p�\���_ˌ�T�jr���ť�pn�IYezR���������q�yg�H�ʃ2jlE�_m���V~;��ũ�C���^	��l��Wk�#�Sw�q&�4Ӯ,��(	@Z�.m5��-�Ω��m+i��QSۏΚ�V�}yL��{Wx;�KAU���M�=�E�w�#��|���3�U8�\�@��=Kom[cn�Ԡ��Glom`iCsf�St�5s��5Y�7����f�,�7��Ψ���DJ��)�x��ջ|i���\��#��nyH���a�T��2��X�f�����A[���Q�!ݘ�V3GQM�x�3��s��C��v�Rb�jCQ<R�Yn�`�%�����ZpW,��\���B�s*w�KW����2os'�ñ_�<#�m&�E"罸8��'[�������1�_��V�ǘ�7���'��1+ϸ��vޅ���y]?���K3z_O[D���cn�m#d��xF.�-���w�����/_M�sj#.�Q@�� �MjcF\d��Y�l6	R �)4g���c|B�ʍb�^mmv�j�%r�.�&;5��P��z�K������!|H#4K�ܤ _v�c�)R�v,�џ�q����{o�s�k�ZIR��mߟ���*L����Mt��$�똲7��#^��*��Y:�3����}����T)w
sk�.^�蠔%|����0��:;.z���a�+=�38Z��y%A�L��wv8L�JA]nc��^���^�9�ۦ5����)C�v�VK�o��"�����_^�(u붖��pM^5K��g�IqMY��*:�ϷX�f�_GAY��	`֘�����a�=}�Z��/
H�m�6�6�I�p�2��d�v-�����4_�7�9�t�5�6�g�`����n*u���Ͳ�T�z��\{B�-���-s� ����M�p-�Q�۽�b�W�����swk*���M��)�[Pus��vac�k�0�q�ՐoCwyz��ܡ�b���U�1M� �>��̳*��{S9�۸]���.�J�s��v�|���kk�m�8{�Q#	I�	$�b���G�E}���в��_�|�sCNW͕8��kj*е��e ���e�w� �A��(�E/z�
������)h�QI$ ��"+ ���>��y�4��9��8��*
H �0���EnNo�_~�}����� :NjC����@�<sq���P|�3��I(�/:�}�gI�龮u�lb�a��l�<�ş6�\�:
��0��xqyp�4�����t��Hl��QQ}�!%�6���k���}����������!��iڡ�~_@�����ʿ�u|;HC4��L�?=����[콫0�yC�b��4�h@
�Vyp�7,�ß��A�?}�Bѥ�3���\�PRZ QPYT3`� wDE�w�	3-�g�Ե���4O��741ܦ�9A���j���c����q4'-��j<M7op>:��'�<��z�XwYQQngu�z)�N�~��lO���M��^]u�r�QM����'7JxsW�5���QQy�P�<�g ��ܯ*���\��c���N/<T^��(�����EꞬ�d>J�Y:�`69�#��62 8,� ��\�a�X�����@@��s�0�_��>� �,��4�(��M7e�2p�v���c$����f���hs���l���
*/w�\��t���ܥ���n��y������y�����}����#��/����ࢢ�Z��� ���~T����=X?���2��k�M����A�%ȑ�zy4X!�V�֙���O�pG�ٯ��4��U�0� �l�-��T[���P�.nn�����9���gnm��e��k�S �J;�����'!��Ox�����3����[�X���c���?���0�^z���XN�G~d����"�(H ѡ 