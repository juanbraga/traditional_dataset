BZh91AY&SY�8�  ߀Px����߰����`?� r$�( �$�S�mM�M=H�̑� j6�d����&�����24hɦ 1�	���dɓ#	�i�F& �*~�O�<�� 4hd�   sbh0�2d��`�i���!�H� ��Bh�)�M=����i����*1"B�	X	?��� ���b�w��k��M�wL �Gc�$�U��_�߳��tw "1L���Z���FN�qjt��#�Ln� �H�@�6*N>y��9�ͨ&bl���!��ը������M�d�H+IIz�����]�	��z���O]�K�����y�]�t��t�g>���BU�:�t��\��#$C̔m���TՁ�C�"����]sũyj[Y�S�܏��8d��Q$A+ZP��hW�iwש`�)�o3&J:�0*����b�5XԴf��I�GLcL0*��.[�'�m�Ze��E�V[�R�6EԴ�m�ګZ�\;��F�0�2��T��������0w�hU�0���M�',�gu���a�)-k�ubl9��l��kK���*��H3������}:♝�D�g���qd���6ɡ��Hʼ�?����͚ˣ)`�H�{�dn��Q�ʝ�CV�K9�%����1$	>2I`�8.��R萻<s*P�+9U�mT�P;�sW2!�J�di>�DK��h$8k������^*�9��3$�m73���_�����M<�6���'����g�<|u쬤����,��i�]��JqX�
�|�r��gRc����;̏�#��@@���?�p��~ޖbKq��
ކ����P�^�k:�Q�3=��R�[�Mc�����x�K�� �A�1�>�Qc��M��B�	�e�U����Ika�(�zg�&�|��T��A��~��Y�`�X�",7�I'.�D(S�F~%�<fI�=�8�Yp
�;��A���6���մ�ENtę����q�F��f��R�f �%��;���[�;��$z.P��J��ݙ�j7�ss�9��xeM���
�km1�ˠ�����R���T�IB� i�yO0��Z:��ja�{��(	��S���J�R���4L���\�iAK6I8L�B�� �6+*�+$�M@J�&�zJ	 �cM�~"?��6� ���*.��9jRuƲ�)C�D��sڜRW&{�`�V�hu]�1Zlb=��D��$�hy�hiB�"��5x�e�4��fI��1�q٨�)���g9m����lI]�acQ|�1��=�
��� X�O��7L��5�5Y`]}�<���۳�4i4͆�d�{�
��)Eʣ3nA��@,L˘ȣ6��0d2dj������)�y���