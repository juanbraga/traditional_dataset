BZh91AY&SY}$d� �_�py����߰����`�z����� n���`h��F�d   4  �56�)*x�       ���)��i 4     MD�DoQ�M3Mj ��9�FC&h�`�4h�2d`  �! $�4�i53)�L4M4 �5� � �B� %P���V�I1$y�?ތ���@2�
0��±(�j$
�B=�)�3f�9���y�����3aH

�T����h��DDY-%��!�a) ����,��|Ϩ��݋];���PТs���g��4�WXʪ���/���SH�"L�H8EU�a4�tȱN�Bvd���z ��U|��TK�n����ju7腌��=S�ټ�t�4b]�;�4�b�Q-���gg��hS�գ��u��.�@g�-��'���E�F<w�w9�>�(�s���Wv� ���6���b�`y.d�<%�(d��
0M��h0m\*'<X�`(b 00�	��&� 	eu��6ۜZ�ƚ&����Fh��	�H/H��襕yj逑7x�39҇�`�`����*���!�ƹu$�*���6�X(��-��Mk4�]tnE��57Yw�k6ɛ&�Rr���]U]�}�+������;l�Xӕۚ@NX����0��!�kn�p!lZ(()Rk����1������縉`ڌMi`�!�J(S30E&h��D"C�-B�*�.V�ɋ.��]�b&Z+�<$=��F���B+�̨P����O���l+�Z�F�9��j� ݙ�;V]P�+����戁��n��q�2�6I4�X�\^
�h�w��P���0*���'8���g��n���K�}�v�S���ʩL�:K�%�Q�{Lë�kk�0ʣo���B��QEN6,F�1��sH_b�}��,��NԬ�!{�ma>p�p�!��F뫤��V"���P��JQ�2�E�!��0B$d:��R��-��I�+7��|8B����8*ER�v���y���� :R6� �猅fXq��/�ٜ��q��<�؟)5�J���HʋX��蚊�����C֦�K�T��2;���6v�0���P�SPoΒއ���8@��k<]�� ����	~]��śo�bjK-��R�+�B��8�3���T��/��A!Js0��xm،$$��0@�/)�N�*�J2F/�H��j⋂J��!�:�Kn)Q�jܐϗ�[)Dxx���	pa�1*��d�NR�T&�A�%`�l(e�&Bǥ.*^=L�ʏ��bUp�A	�`^�n�0`���o��n��lu%�q;�r��ĪwN�%�z6�Y�AQ����Dؔ�����/M�|�����I���݃Eۘ�	���`k7U׼����P�4ȩER�[�A!Qu�2a��E�~�Ls���%�� 7�4H:��P#x(��`y�4Jk �^��HJ�$izD����AlU�Ls����I#ID2�^X�HA�ń�ǻ9�PC�Yd��(ġ�Vx�C*)R�䈥�օbJ�
\�D�i���Q��FC�5�� ��rB�W�!n�$��ю�����FI7c��S k��R��])2F�C���+�62�N��v���F7e�:���(N�s�|A
2��Z�����c>Q6�W4�b=w��CtY%'��a[%*�c9��n�jL9���y͓1P����9j�[0\MW�Ō2�AF�Mf)���M)�	
���^��a~�f�҉��J�	)�e�&nD��^�%R��<�ߗ�]�s:�QXTb����d��O��u�1����FP�ϙ;5)��.�p� �H��