BZh91AY&SY��iD ~_�Px����߰����P�9��Q�ƊQ��$�4�Mh���z�ʛI����Si���1Jh �     �)4� 4   �4 9�#� �&���0F&(�!FOQ螛E�i� �@���@+h�QQ(�*�Ft���A��Y�/��B�i���(7b_	l
D/�H��1�u�i�G�	�� p`�>8��t�v�-^�0��3��1�7N�T�P��(��xv*�ҵ�k? ��"m���0��g*����-�R���|��I����i@�O.P��Q�א�����:v;쾪�|��n���GsoVvqt͍�1|+!8E��n����Vk8w�j]�um�l�(�P�ִ8�ԐaD����0��ڋL]�
m�(HB�e���T�Q7ܩ1��,"�Ab��$(�T:X�<��WUb����@���;C<�I�GK��˧�o�7��e*J��l��SX�"P�A�WB:		Vz�G�9d+M@�4��K-M)C��YVPK��k�4i��K��U
�
N������5�Y& Ԛm���X  7� ThP��O^�T5m�Y�_v�SV�R�&	F\�C`�?JE!�?� �s(�kt@B���1����u��aT[�`��@��c�.�'W��T�=zo�9K�����?�����������~u����$ ^���+�B@�⿤&�]Uw|��XQ�u���Y�P��:�I!y�=X�	ϦAWj`� ��I��wN�ӝj�KA�����	��_��;^}g����G��c��tmf����ނ8	���<{bL��6~ �r�*NZj���:t���!�����.$�E���S�4e���h8����iX�KH�p&'>�[/LL�a���~8�R��I�1 ��}bB=ˆh�зkNv��6��P��s�ѶD�8�e�G:ѡ�4�ea1��Vi5�j�D̹��j�V�#y�+50̘l&��}1M����B�637P���'� �H]����r1c�T�7���9q���E���b�&�+( $7�Ž\ā�Z!�5	�=�
j��������·���3���Dh�	���(��~�;"�����v��XҔ}Q���A�������e�v#Ұ��6�=��`�X��&�aɣzK��sv��k<��58HNO��O�d�-��|(^��Ƣ�Ԙb"m�bF(|q����+�M��*�x:S�(�iP�|�U-��a"%-h	
L M`�&��蹇(�ҥw"�N��F�`�� �ND�L�p��/��pl�d��;m�*��^�th3���@�fGq�F�'^س\��� �wl���)��3J 