BZh91AY&SYڍ� ��_�py����߰����`��|�7
T�ahQ `�	U]�         1��Nw��    ���4�v�I���b&`(�݇\@4PJN�R���(��J�@ʌ�F��F�� ��lf��h(H��b�@F����SY5��4 
� Ҫ�����)Q�f�
Wl�h�M0�m�(��4�c+  0im���P��J!1M"Xl
���1� ;� �ĒT0�T��	�����l�Ս��Qm��� wR��@�� %ID�44d  �� T���%USF �     dɦ�L����0Fh� 3*�EJ�    `0F � d@ɥ<i5=0)�f���$�A
R�eM   �� 4�hݖ2�)ײs�%�ұ�A[l��Ȋ ��Q���)!UqS�A�d ������u?��`� ?t�@�!Y���CUV��5$��		PaB�B�fέ�I���쮜�����aT!�RH �� T,���B��A@��&0�@	VE�!R$$X ,�R@��Ld �@&� ���HAH�
�* � *��$b g���C���C��ϻT�?�/�M/ߐaJ���vE�����kUk3��-�$bı�J�Ј�=���Ŕ��V�6]�x7+^�.�\�X�uz��Y�j^?淺��YOW#����rc�u�^'�"����H����v�C�lHYL%FHBܧt�ˉ�ZY�\rV��ل�%�IS/.�.��)V��F'���[M�fm��B�ba�j�,�Pb��%bmM3���˶d̙�CX�:a��ٳ�M۠��Sm�c>�2��M����������F>��)�"��<"�E�k$V8��u�{vIOs �v-��w��Kre�BQ�� c����P6�m�/�"��L�R&�J�{4��+ˋ^퍻�q�P�()�Wr��B�G0��K����Dn�1 A2��e+_�	�y���V�3��C%ё;SMV��3�J ]3�j�K�[s@�]�ٲ����W����;J�'%�ͻ�"մ.diZ:��[�85
ur����� ˧.V�7@���c��wy�R��^�������	Yy��s�O9��̫��xh��Z��\1P����_"f[T�	"�D��Y�d㳻t
L�9�;�-�sD���������~Q�`�`q��I�I���DU��AE���G�Qh���Tb�P�Qb�ݾ����"4�y�7(ۺQ�k���7a�AU|p�(K!�1!d���'Q`�[&Pٰi����D? �B�5�u��/������v���/i�ע#�-0%-��idՕ�3.�LE�q���w��-1��[�$��42]�?T�.' [��B sN	kh�3D�not�2^���!���T�d�:iQy�q�s�����-��2ʶ�+���dR�,L��d]<A���p ��1��rsV�� �伫0L��0# (�8.%��ˤ�K��*[շ�1"Zݦ��ͽ��IB�y�?;	MZ���/�{�:Y��9���Cv�)PyWlT�Mږ2�/u{�P�P��5��]���Q	��V�5F)�F�U���;0�V��k��V���J���mR��
���g�.��v���6e<��1�y�⇬��M�w�J�k)fe޹uu烺y�t�9�C��x��'����5��E�L��6��+����W�0�ѵh�/�8r���Q/O�Vc�G� �2/� �&Zr��-�pQ�IU7L�he8"E��N��c(](
�	qv� 1RQ"�aQR�y�3a%%5.m7��dm��-��a��������`JF[k$�f�1cn���Ʃ�h��e:��ևt�ufe��S�W�Y�1
�l� d͖`�$�G)��SX��� 衑F�Dm@����TQ��I?;��.���j��d��tGX�	X,̬@��oM���tsVj{c�$��kV��6:7,P�jr��퍠M�y���CaqMDۥ��B)+������-�if��ɛZ�L��&��N�A��]d6n��"U�Q$�..��I�"���M�d@4�'(�bB�c�$�g�m$v�$4dG���f%c&I �i�KHL��U�͉,�0e��e�Q����,���z���l�Ba�����f�x!Ëd��Vƅ4A�4e��ɹi�[т���h�BCp�@Ƙ���K)D��2���.�V'b"����v�	�c��h�����e����~��?R]~�Pk��^��y�ɮS[�-q�ֲ�7
0�6����i���P�`T̎��&ۂ�sm)SiT	�.ՃMvƺ�f�6;i�=�������q	[pRR]�"�ʉ�n
C��']�M`�3k2� �E�t.�R$��.�K���M��Q�m+�hb������k�x��;k��9�m5�m&�3 Ѷ��˭�3�bd
m�v����̺˻S,��0�h�(Lh�˃��2�������J٦���Ӷ֒�f.��.�)N��F��Z33��47b�]f3��D&�K*��-эt�D��[,�[��f��aI�	k��ى�!f	U�4w)v��(��Z8�Ĵ��L�ͱ�)��]e+����ZS;��pK�.��H�(݂\ƙ1�!l�nL�u�7�Z�^l6�[\�Z�st��h�	�L$�6Y��m�j�#��)�*j`݋���ZGm�2:벺.7u+n�;X��].��c��붚�7�fmd,֒�K�H�f�т��*��Ė90��[򆖶=�����Vkv)�eJ�Ҧ��d[��*�v��# ��i�:�[���62R����a��u�QFې�%4�".��B��XX�Z;��(�MSYl�]5˩nh�1;XV)�s�S�C�P�$���F,Ĭ������%+�.�LSu����#Bm)6��GMr.��V�MN��R�\��(��� [n�)uI�T����V�tKMv���6��y�i����
cD
�)	mynie���+abX��%��5-͖��iYSu��YM5*n�l�UFѦ�ike� f�&��s����m��t�nyu�ל��hҵ��M(������j�9%ZYc.,e�k��W�P#A[-Sd��1T��\�uUXM��ҳ%���G�7;h�Z��0�W��ŕ�Ґ�΋��K�k���U�m,�n�悎)B(�d��YV��]�!e��u�L��ћD�#��ZR��h���,Q���Ͷca��١-cmc]RWY[�J[-�]���m���ܢ�-e���6t��FU�`.��5m5%nV�"񍳻/n�,v�-a.u�n ��B�A �]n"����GnԳ
[M�u�v&�B���H�i�/Q�%�!,me�"a3+T#n����8�M͙Ve4��v��6۞M�5�Gmu#+�C]�U����Vz���FYn�d��v����6�\l���B;f� 9��1����=��7�����ƅ��L�[�K�u���q+�mF�S%
f��Yqn��H��X�z)[����w� �5H�DP[i�����y}����1H���!<Am���EK�Dr�L ]p�� W��ݰ$X?��	��$�m�
�i�CL��)&�'���?��<q$�HC�!���@��L�:�Ci&$��0�L�8ɏu����V�s �m=������&�l:�9C=��$3tS�����W�.���鈅�伵�DC,�ޚ����έy��nSv5X�T��;M7�y-�9�s��yi�����N�����ī�均�f���)��ʊ]iʱ��V�r��'�.5�$LK-L�ٜ֚lk���Ys5���B��5��C23���n��M������d	���;U.�b�"�L��{�Kw7au���[�-�O�ӳM����g�����PV""!�s��4������;��o[E=��v���o�Y=��� �#���Ю���D�V�V��Qr���e�l��.�x^Ib�n Skt�jٌ�.���i\�5�SM��6bh6gZN@�Z!Ku�[`R6 �B!eҥ&�vu�t��m!+���q�Xճi�x��MKK�+2���)hm�.�%�l��m�)���(-ű�gM���J�kR7�Ү+ uqQz�M��-lR̝n6{ld�8.ɝ��L�G&�:䅣��!
%��u�bS���զ3b�L���e��Pu@Kэӣ-�fTr��kaC�쐄9;ܗך���uΉ���h��@!eՌ�1tjņ����fͨ�u�Ѹ�LT
�YBɬ��r䫗0��7�~�$� �H
�a'�h?F%`
���F�`@yܒHghC=̪����z�
����h��X�#"�TX1AQDQTUAX��V(�&���5J��(*���1�U����E���* �"�<�n��*�""��EEb �V��b"�PF$b�*� ���QEQ�J¨*�o[��"��ET*�V(*�� �wlQT��X�X��EEDV)���Y�X�#��EAVDEDX���7j*�_l�}J#8�������DE^P���U�-¦YQ�b��V=j�*�Q���/2�������5TV1#DV,�A���aE�R�:!]�U��E��1��"*#��;jLlb+��*XS����YYPO�"���B���4AT�H���#�Ԭ�b���H�ը�`�kv�/8,EU��U*���SM�(�(�"(���X��X�UO���H�֪��`�6��USv�7j,EEV(���s�s�h� ��7,�V,���M}绦�Q���C�[j���S�UU�U�(�~��v͢*1F"�*��ȣ���b��DX������	�[�c#����{N�7�W�u�Vݚ�v]�y��|�q�(".v�DQ�+�ʩ��֢��#�钴~癤b*��[J���W9���ALJ�T֊�.e��&"������
�(Ǿ9����移�=�ͷX�X%���:qh�
����� $O��2����E�Ԫȥij�,Tc�E��ZQ7��)����洧YE����_|f�(��.5E�FбW�Y0`x�E�YX�h��n�<͌XǟPď�U�,Xow�W�i����E�����A�Z�DUP�Z؞�0QF�1�EE�*.�Hb��W�2��J�(����xq���`�﷚֠�LX�fQ��5��׎�X8ب�}�s�����PG-g�Lj_�*���_'ɮ��MK��D�����_�KՀ�ԋ�Tݢ(�g���q3/<���a�m��E�FT4����O�<�˲qA�QN�r/{�s���Ԩ]fOig�AD�\9j�J�Qz�ϛa�8b�{��I�>ύ1F�^2������U@-B }�Z|��{=�9AIX�&�7�|+w�y>F33�<���"��Q\O~;χg\�N�j�����W�D{|pY�S7s��M��ˉY�9�b���[�uz�^�*�Koޗ�n�b	xY�ᚰ�1���"��Ĵ���hQM�Эkm7n�3<��X�"S͞�u�㥺�����aC��e�k��,��m��KQf��E�v�;s
�ϾѾ։�W"���f��{��c�U��7,+���{5�_-1R��Y�YKue�ˉ�S�xq�E��\�c^�4�����V
�0=o)�Wm��yq�Ugm��V�O|��b!�1�̾��_n}�J��\�C�ǽt� $u��)x������˷5�")�*��o�Ͻǒ/R��>pR �wp/Z`���/.�k���Z��N|�@�&N��8�Z����G/Ϛk��{����E���=֧-5�bĶ�Bzn˘�� �lR�Q��HE��
��Z/��T��y��~���u��c/y��:ɾ�B��k�u�
*��f;��9�d�{�Ň��P^�fӜ���7������ SP`�1��c7�/{�q<i�b���>�ںO���O����e�wZuN�b�P?P(B�I��2��	�����}?,aU�#�&	Q0	A�)����u3e�630Lk.���K4���̫��űv��Y���c:�����fb̍�%�ֵ��~!橈)��Q���+\��1?{'7{r4}EL�_D��������"�x�8�fP�P�m}.i�0�T� ��7���X��>�_,�%q��7 �z���]���u]�.1��,��P EAG��q�\=�F�l���lo�Y��C����E}�(��r�'����ϟR�Q�5v;&{����/�,��d����K��g�!/�:&�+���o�����{���}�mHO���I��� �@8Ã�*��Ěd!�l�CĜ`��I�,�H��� �#|G�j$�c��C���#Z���L@,("=7�F���ø�!��`�:R�HF�6��Q���=N꺤��7ۙF6.����56��ۆ�S����MD�P�
��;�5���]�z��K�]Y��t+��.={��N&��7Mz���}]~����|�A .ܹKj�J*�P�a� �.ea1W���iaqB�]Pf4E���������aB��1Bb#�9!�x����!��;��;2ɋ0�ޙBL;6W�SP�̥�h�P�20�l;�>=QB64��ɱ!V��C���"L��rU]�8Cﶌ}�7����>��t�� k������6�6& ��9QZ\?�������_GvʹH�& ����7&$[?DX�`��x��Ɯ�e��X�" 0`��W�穊�r
��~��������-Dd}&��c��$j���8��_1c	�ˢ*WY���Ӂ�W*V��)H"d�"0A��a}�i�}�;��W8GBh�{?,�>|�����aA��oG�!yN��v�����f�R#���a�,D�g�
�����N� ەU垨���~�I���r��ݙ�&��>�!�Lu=q�pxZ���X�qq�,�"�SN�zw?U�?+c�g��nsƢv�۸k��"�V�%\J$�,0Sn"��7�c�d�&�m ��ҖbWB-��Y�Ҳ�1Bh�4+Ơ�R���
,G�ԭ�[-7 ���J0�&�Awiē�b8`+D	����ڎ����쑥��u(�
$�k�R!Z�䘫ނ�~��˄D�y?`���|�&0c���:�C��݆ÜQ� �*aD��c���(F,��!B8[aD�#�&�h���߆�+%'� �Z6[X2` E�a�#D*��!e�w����V�;~�f��W��Y*+�^%]��J�Q��4�>�* ���A�`
�j�X��&c#L���q��
4@��mM��| �l��#8��%��"�RlCڴP
�]{yU�SaV3[�$W=@38 �2!�%��p	m��p����H� ��K�7h�E���hn�� ��"�:�`��LL"F��و��P�~¶�MgD}���+��"ei��Ф\eq*�i�a$�]�ִ����ҡ��睮��]�4�s���F�[���Ӷ1�4�(���Uj�v�XW,�ɠ��n��m�@X�V����i����3��Z\m�Ux���nQ%u󘁾����Ccm���hV��u���lT6�c#J�6)�6�����y�9��
�	�p�7�֭�3����ˎ��" �d���4�,  ���"d�$@#��]~�1�����w��������bCx2�0,�cF(GIp	$ ������Rb�M�4س��"p0`hUp�Lpe�(��,���F$   | zډ'&m���q6�o3�S��m+�TNRǏ_33�F�#�MyӋ����;�a�,�"�� B��#�h"<�����9�??.��z�E���v��0�I<H�g� B� �9��pX(�{�y�����q�)���ֺ�W-^�߹�5��C�Οj��s��9R�mP����e�39�p|� ���s" ��<\6��_�/U=M���SEwk�����_��z�p�P����_p��m����I�����H�%1����i���GJL�!G���<��DY�  �s��i�gߙ�P�v�zՈ���{��*/���l�r�S�� ��	����8b����b'|�(q$�!|�F &�[1z�ƈ�d@�L�s&�vX�2�P"@�����8|� ;sV�m,���=����x�\TW�`��\>�2:O�f<�PX1L  	�`f���N�X-8�Ti��R�2�ZB�o���Pӄ[�5��v�I�Ląѡ��֤@s��͕�HЗd`cQ��L�;`a��1vL�kY�k8|���o��8r��9��m��$Ṅ8�ǉ�醾  0���M��R���~4����z��}�b�b Q�M����1�C�a@��\����`�Ծ���^>��� ����ΡAXb��ރ0��ۭ��xj̉!$�?d��  DY2`ňЄ�o�,0Fe��Ɋ��LX��ds��w��5=|ʡ�4m�nS	��� ����c�+D��l��Ӫk<Sl_�XT��4��2���&�/�������+���.�X�, "��#�c��剘��(��������PҫP�}j�Tn��T�� W��� ��4�T"`i�"Dl�̦+��:ï�;��v��]�Ev<��wFo����M%A������ɖ��.�{�.l8�����\��m���sp�?/a�F �Y:b.���m��7h�cd��O^��ѽ�tg�|�В"bD6 �r��O�����/sS��L1���4h��@DN�&"����9΄V�[�&�$�;�|����TmX��g�)Q�yQQ���(B_ ɀ:���Y2������
� ���"4B��7�'�$�1ǂ}U��uP����q� �C��i���@'�eQ� �5'ýJ8�"�q���� �W��z�6�4���DX�Dԯ�;�oĉ �(�Ǉ�pt�g��c� �J>�0��4�|���6�����yt�������5�m��3.*�0�e�����@��`A�8a)��~��M@�F����ykԪ����ek��8��6=n����Bus�� �@�+M�k�;O�>B	��0*�ЄF��""�	�Y1 � aRc���x`#��,�χ�w���q)���#.]�r|n�����t,�RV�d.�r'�"` d���́�D� }��h��f���ﴻ�nĩ�&?�����A!�Y��#���}b)+4S�������ˉ�Js�1'�L��h5� ��%���Z�#^���*,�%:�G�r@���B�A�qx����Vh�}V�s�+f��Ϫw�� �u1z9�6�V�`�s,��&h�q-&R���h�Z�:H�fX�u���'�r�+03"�w���}��x��-���V+!� 򊇬���X��[��~�P����S���Jz��@�ip!BB)xm��D?�\
��D���V]wdI�H��ˢ�1]��vH�V4��\��oׂ��8��-�(,�(p�)8�@O��Y��f��uS'�f���U������w�(U�A�>�l6�G��D(
2�L%Wq[��̛�q�0q���㜆�����-E"w ]6P��ĳ���O2���R�FI���	A����M�I��v�OzfA�
���E�[}��\%�}@]��8�M��1H�٭s+J
����}��;O�G
�G�&���C�# D�8t��	�o���0h�I¢��ʠJp=�s5!�Ё.����10J�v ]7s8bA�5�힩7�-K���ٳ����ۂ"bI�Fۜ���i{fDW�<��Ѵ��+~ݐx^̝�{�~�(!�*G�f�h�Gm��{3�&8�Z���֛qFy�٫��ZTGb̙;6�����NP76�N��}y�����3^(n�E����Nw]�:W��8P�i2�n6c�2�1�&&c�^��2��zs�/�GĘԈ�ũ+u1ә�ɴ)p?���\pH��+�V��%C&ǚ��+��e�<�>�j �HoA���'gEΩRL��r�3@���-����4Rx(�:F	�5#��R�۴ƫF#�����0ზ\��	hڳ�9��RWH�V�)/[��dd◝
�8�j���q1�Л��3�Fƣ���%Ⱥ�@���;�+t�ib�Z#�7w�i5�-�$��z����0.����[{��]��x��
g�ob*��;x��E�ۛێ
�.;��店oE����>o}�m��=~yC�4���k`ѷ6�%ip�m�k��I�[���7�b�MĶ8�lK`�V�R�A+k�`�v�ݦ�$m���c5*Z�J�6�vۆ�֣�^F))	�V;e��1E�,tq\R�fe��m��+�ض�R��*�����γZ��%TLā�(ӆ��,�i�J��ė�̶��eP��Փ%����A�!KR�Ȉ�\f�$+��VR6�L[\���nF���㣛���U���.m[.��g"�����N�����S߽���-���Q��&�qF�n�:�E*�ܔ����#�c�$3� F	���K�9.fF�A�߯��~�͞
[��5b�O���>�Q�-z������}�<.u��@]�� �כKҾ�}+��na����̀,Z����9�� r�ഭe�:�V�D��
��Gtp���H��8H8(�i���F����;;�Sc�2\&Lt�(��e-ˍ5����Q]�����gawv(�e=eО��}&4Ӳ�����%*�?(^@[h�Ȳ����xV���˵�!R��+Rk\!�qb�������k���b}~}�����Z#4�HŪ���_����ڼ��TH�D?��Cnh	,d,4��[q�[�{�r�n؃�Zׅz�ۘ��A���P���a��`'8YF�x���e���i)[���*	��%3ҫ�Wh�\�h)V��?t��V�C?�����~���$��L�j䫔�5Ң��U^v����O޸�P(R@��< �p55�$�W���'ד�t�;1=_PJg�}�ݨ��Xzc��8��u��ןb�/�TbQ��N6�0��s#B~��uy
���m�c�~{�VϾ�����5F���_V�D!ٗ&m(lR��Y�A&��f��S(K
�Ә����B���@�l�� F�9�^P��0���܂���,T�`��S����L[�s&6��K�wQ#˔>z.ȼ��%z����К�20��B�e"��m���l�b�"5
�v�f�rlA�T6�eu�isGg5F���m��h͝Րۃ�u�3t��0�")�y޹e�5.�����H���P��C=N�x����T!���ډ�^�K��딕�+�=M@�+��h?N�f �!.�t�nV�>;Y���|�)5;�?!C��B����$�
mCd\�dq��S�ə���_X��}��P>��Pm���qս��Z77TfUV�
W��p�0kKqC�(��q�^���q���K.MҗDr��^?����pI���*{��6z��W��&u�+?!I��k�|˩�+��z)�h��fLJ%Ĺ�? �-��U�.Y5::2;0�����^Hʴ���B�,9�|=�M�lR:v�xv�g�\�Q�/�\�%h#���0̂���f��r�g��Q�ԛ�bl;F��ɤ������cd�.�!E��D�(6�7�	��߼����(y3K�34��^ݬBP��˴D�h*�w�NUP�#�P��V�]�᭞�!KeA�mѼUS�2"cBq�DB���aۖ,u�}g��q��u9��1l��M2t��ВZ\M�M�Zj}��V}�z���j��]�ȃ��b�.�Z�2(���1`�>5�5@�̇wW$�2mz��^��Lh���[�yw3���B0�S��Q1��ܞ����>��כR*pW�gr[�a�Qq2�N�����9˘Ѫ�j�k�H�F��K��b紸2\�u�R�	f�Қ�%��Й�݋,E�R��Rǳ6Ηe\[�Ռ�Z�N �ۺ��9���->6z�P�=����� :<�E��sYg�~Yy҆R��[���|��`����s�I9|a�D�9�$wd�ਘ���{;ͼ����d�HE��yP(.�e�0�6�);�w}+f��F���4�2Qwޝs�X�߅��v5��Z�J�Eoff�g?o�;���T�u�G���q�M�D��#I��zp�~��E/Q�����|�l{�	ޣO�����]޷	������E�\Il"W䟀�@�iF���4��ZY��X��^s���B�-��"������_4f�Vb^xQ��96a��v���;Z���-�- �Bη+F�j��fN�}^�Y�TR�YJjR�k�����p�$��V��P�[�Ԝa��f<;XUh{�zf#uws!�nc�f.ݻ&�qow)�[{���̅�T���]<!�{[��.��ٙΦZ��	ݸ#P�%>��7y�CP�yB"��^&R٭��v�GJ�2]�`w�n	��@�����q��v��*e�ډ��=#b�b1(ɡ1��Q�C6���8���ǻ��:n����<�����T��kf&�E����a�)�R-��׼r�X�-������?|�c�H�f��4=L��%~����s �N'��my��0��g�ڿ��5cD�m��]F�����+��N����w�Z�T�0~(ـKl&Ze�9�g;1R�����6�K=�(0��4�Ҵ]_��TI$��P1�MW����9$W�Q9p�Q,�^��YQ���%���^�m�hw,�3[�b-cdp�7��F�y̽T�j��S?'���9��@Jk�+WR�$��F�٘6PC2��9��L��G���lu�N�m��a�f&�����Z%�X��-ǯ�}�UM������m~tc��S�;���3"��:�;�4��G���V��VP�0x9Fj�����]������.�ň̶��쩑�P����
��<�(���b�I� ��FA����B �wnb�~=j#o{Z�}�`&�r��n��=]5�a� s����l��w3��np�U�E��ъo��=���ѾU7=���ظΤ�X0���ڌʂ�kÖ5�rn*EԀ �m�گ�s��dA��	��	�D�dC
�U�����k�]�P�D��s�e7�4.���/.���=����������RgSrgd�.�z~������j��H��R��ث��׹����tcqd��L���U=o�&=z5������Ш\�s&��D��r�tsʝ�n\�����"�S�J}���^�\5����wܓ��(J��b[���,��{��V#�L<],�?y$�vwN�Pcl�Vկ)����*��rvH�ۇ��"��*��4����ߟ/愾��~u�talf�T�rq@cT)��R15���ӄ؉zOP�
��N//�:��Ngǎ^��B�p�;������/Ê�#m�j�Q��/�U��c��1m��:��0A��t���S�=���u��.�h�S��$�!2ɀ�$�66�n����u��kF�&��l�N3̬#��GG��&�g[Z�	�G6�mu+M���.�I"g<)LR���/N�>̿"X^+m�U0���@���RG�&R��O�ʰ�m{�U˄��J�Ƒ�$ך��X"=�!<�@�w��a��C8A���R	�
P[�Y`q��S�1���=�V���@�Ug����]B���`�Ҍ�T�*ٷ+��R��ڞ��Y�ĲW�@�/���dV/CJ�n_J�r_s�jb���5�b�d=NqK �۸P\�����ȹ-@A�7��d%�Wd�T�引s�z�N���8z65�A��P���Ƭ��ԑ�u�Y�`�fT��x�oJ�����&��M5���1_f4f�*Y�v�)Q(y<�=��� �o�ӄs�velp�=�"z�[&��̼Dm�;07�_i�� ��b ��;C����AĘ�W�ۜ��+͕�9'��r%97&���k���D�>�{��Sw��k7&32���"G����=�S��u�T��� o�d��i�߶��S�����i?��������<�I�d�ipT���)��1מ;�N5,��c�7Scu�  �"�=��5��W�A��kۙ��ξ�a��s�B���$U��]�W�΢��z�-`ݟ��:�Z��|=�B�ރ�w~�ٛ,	�ԅ��̒b*$�,���r�4�g��>����$��A
z77�+�^?�X��Y���ݙf�d_2�
1��P�����M�"C�������
��v�']5��'oD:��r*�R�DX(=t��FF��]��sU�u�I��RwɖK�9t�b�����8����	ܠ��,N�2��X��%I�E���� ���`)�V�ϟ%o�jY�k�鵯�%��]���3	]����0ƛ^4�M�qn1n����u�Q���5X[e�U�a�r��ܙ�)�c�����Z둗k3J���4+.�������XD3�"C]u^�kz�]b�c0���Il��6j�͖hm������4ieDX��ɯhWs��-�v����7LCs��P�V�����b�ҕ��n�h����u��#��ˉ�4h�5�*��bqk!-�g1�#5v��x�YtՍ�#��] ��Śt�����}�9`�]P�\�S�����s����Aw���mr.�vrlTG&��E�WnX��J��εU�g���3���ud����{���ILX�2v��+>�"Vf��>�0L����w=�? ���dR7�� K ��;��$Ir�Q��.����t���[��ˤm�֝��wۤ4p��^� (*�7���Z4[J�`��l���>�K�Ђ�m�f�r��r�xԳ�n\��؋)#�
�"J6A�FƀZ7���V���#/1�ȿ�o`�D6ߩn�F�mt�V�åN���a����Thj����j���
l	?�$�����Puk-e4nZ�Y�IaVY1������Kv�e�lT�9��ީ�c]��7n�^5��٭VRB��3@�x�;Dܬ54i��������i�}����r5��;
�p�,�E�L��N�F��&�ם��Ty��!������S;��7������4�]	�լN�������7~�|��U�x��h�I�'�,97qz�-+����^��~&*{7��� ^򍜅��)Q%�}G��9��)'
 ��Bm�.+��FK岁0
����:��jwo����Ø��B�;���4:"�с�];�G�&� �Z U��7����5��W�o�X�AX��y�V�|wF�d]otڨ�y"�GJ�b������}�OozSL:[�eq]��q"�b(�e�ʩ1iV���q�`VW��u�\0���5|��v�3E�p&ﴶv��4�슸��`\5�ŧ}�@�6'l/x�ĝ��z){
���X�pz"����R�����,���Z ��Y&��臭�^fO�1×o�=��{�Rbw�AP7�A��0M�W?���{���+���@������Nut��uFf��E�V'�ұ��B�v����⷟�/&\:�v�l��	ݩ$ظqIԥ\�>+����0Q��Z���Z:�E(;y=�1O�5#Ĉ�t6���L��z����i!hٺ�mi_W���:O��8�,��#�AW�W�g��*ap�Νap��6qm�]E���{=,����oi��}�ʍ�����X?��]]�=�Moӻ,:D$��J�V�j&$�8�Pkn~�{�N]�����PCۀUti�WNL>�&�V�9/q���hb�I\�.���;��Q݃�)_}L����������8���{e�Z拼�f:��Y���^��уRʬ<"2,Ǫ�ȣQ%�)�`&�.P�[{OƳ����V�[��k۩����hם��5��D�<�1X���}�G2(��>��8W�3�)x��)m�Z�&�쯼AA=�|b��'�Ѕ�_}��_BִzxEF�a��D�ŏ/� �u�K�[��m��%#�b &�JD�vñV�b��5��vf���ڒU#�b��R��K���޿~������3�W<4:�p��yѲ�����ї�(r��"%t��b��R�w�Ux:��I,Z�RF���!/�fxV�0/�X�7,*�
�-����z=T��z=G+�.�dk���5'�m����&���ɀg(��.Yѫy�tP�d����WKP�g�f�ۇ�ز����o:d����qy�	t�z%������m�a�j�qmCs*�s���=��v��e�3YE�[W^�F��Q��iI&[l�%8�M�6mf-��m���f���_����*�tK��Z3���cWoi�/���<�\��N�b�ɕ��+wS9iF��a�w���� �����tDO琓�'���UQ�7I�4snjs�ꮃ��!.]~�u�O^��P�.q�����Q��Jf�}9*љ;�:u�K�u�u�VJ���kEP��.��1~�mJ6���))-��"r�����73yt�F���V&�?MUSk)���ǹ�lma�"#����<I�m�wL����6���+:��Ğ{����*���0a����a�zΧ��ܾfd�;t�_|�{�[�aS�m��+*8�a�� �}��̚ջ�:i>�菳(i�9�kqM�:�Fl�Ol�Ű#o������N�GU�
���ao�rġ�'������� ��� �!�-�Y����0n�s-0j�:�B˹~o&+x�sShvn7=u���+��&�l}8M�v�V��x��%E��ī��l��y���(
[N��tV�-�!�NW��Y73x��=��=;�{�W	��f��%ʨn�}.�,�e��Y��}ﹽ��[y��3	I���3[Q�γi}Vn���Ku|\y�EX�JZ���y�x���g�{ʎ�2;���=yc��ٿ�V6�r̈́g���R�!�U\/af�|���2�Yx�&��p��9�u��́�d/v4aXҡp�Ipޭm6)��[[���M��͓�)K��1RѮ.�e��4��y]l23s*��_�����������dY&<�Z�&�J-z8�Nةɒ(�w��碽檲t���1Z�ԝ�������'9~�'y���q�P���X����~�9GL7�4ȹ��� Q�	(��e@I�a�}�٬\ݙ^�Fr��F�y�L�>������βѼ���i���o*�}�[B�������옡݋#Kw�݋�>��φ���V�M]�wu^�Io�c4�o�M��_�4�5bWd��C �oA+2')q8v�ٺ~>��!hF�կk���j����W<*����Y�+���-� kQ�uw����֧�t7	��B���>�Ӯ~T}������{�-����e��ԑ��WP���$�eCP��һ���L�vk���]�ɫVu�=��L�r��1�w���qw���,�ۍ/ݺ��I����+�;q������'�{\&<�Ď���WDn�v�r�ݳ�xҋW�Plubp]��`Fh6�~�8x�,�	4K��m���n��EJ��3�;8�?e�������V׶P�@<��B����=K�C|���g��힡b`V�������*a��jґ�X�aZfy�	�ɪ1��"��<u���*�.���.�$�u�.��݆�`��]v�QC[�/Av�9HɋZ]t��au�5�#���?>�=��-�����%��U�eR"�LNlvnܔ���T�og��2��Q[���ʝǌ�ێ�W�&�kH�>�T���JBʞLF��]�Ղ�:����B������D����n�t�w��w/���ia���̜}�v�̧.�s���պY�^Ckk��L4���H�{���3H��tI|����t�q��~O+��(X��U�c�+;�6}Y�"�gcA�ʃK}�R,��B��ZMВ6̳G3s��^��}��u)�9��.˨�Fh�Gl��^�ʋ	]��L�$A� �J7���G��\w/�5�aң�C�\Ȩv-\���=��}�������6���j�����a�����E?J��V;ك³�c�|L{�Ƿ���kp�)t��b��~`fл�͗�|u2��������.�ڬ�܅��6���u0����i��:�/�9ٲݱ�u1�#�޻���ߒ���ٕ`���ߞ~�=��?+�;�"�@e�r�μ0�ܿi��+Yqۺ�+~�tm�n�>�>t/�i�/�pj^�5���J��-�AhNt�WSw|��os��t��Y�nD����d��T�g��џ��/W���͝�razҘKVGiv���1I�L�t>U�a8��=F��	S�����)-z!X�U'�����G�xnqV���d����=8cˆ֌�HJL�̲rV�lL��%�74�e���ob�I�׫3K���u�p�+s	��i\=�ۄ�/^�[� 켒���w�! +�X~�|�x�L�t�Tf��k�Vk�G�k��4Y+�3���q�M^��5
���pt�t[N8i��Ֆ��\4�][*b]����
e.��r*KGD�VLu�m���ڭp��׆��jm)c\���0�svԘcqR\kKv�a�'f�a��lC:�],ڙf֝D� ���j\˘�����X2-�eT�,��L�,5�k�.�L�m8�Y�mmҌ,%J�Z+6��Gm]�KŻ8�֛%��Zk�֗��w�^�\�I61��j�c0�u��*�M�v���b��l��u�g�V�R����6݂�˵a�i �������� ~ҫo�glj�#sq��������8�}~�3J���|7�������b��<�R�C���<���p*�9�B�y��C�,�@P�H������9[y���:��s�z��=ٰx�ů]\�PCU�,Wތڋ']lt{�mVzᭀ:�N��ŷ�+�kZ�p�	ı���f=�J�^v���kޏ�H��؎o�4I2�{�ߐ��t��h�Rf6��<��Ev��'���sY=c# |����LŅ��lr`�{|#�n��ff�%����fevK�a�C��嗮�O�Դ{K�<4\Ƨ��VF5��f{�E��~B ����,��MSH-��U��f&*�
��n�=���l�fM�]m	-���s����6�	�C.k]v�������pc��λ�a�hV�]d�)-�I�кV{��oQW^��ԥ70����L�-��@'�p�5Vʲz�3:����m�Cu�Z!ޅ�p���`�(w�4_�D�L�,��<�z7��*@ټ�
'���/�׍����3��o(l��cR����y9MԚ�/f����6�#��5���`�4�[��P#i�45ob4Mc@�R���F]���@����ZKiG6��u5���~��7��O��ǳ#@Js3�f��bB��pЍc��V�:�4fFouC�R	�����Q,��X3�UThճ��n�WG"CH� (a�I��SB���<�ҩ����ܾ�dl�����V��}�g%�nƹ�X�F�E�չNԹ��[/���A\�ܐ��W����+VGs��.\�m��q�n6�[���v�)R� w]�{�\��]E�9pMC�C�S�$�y�g�˝q����A�r�\{
��;��X'�{+D���u-��>|}�f�T(6|<��/ټ�Y���Y��{3\����l��pb�{����2���O�:�� C��C�IL��Mf�r���$.T���K{J_Ο��D6�V��cZ�]����R�߅�373���iïy�蝓+�c��%�p#���.��`�[ �{\���)��<$g���{
!�Ii��l�-��tT�Q��ͺ]��3����ff�W��P��_�\�Y��lN�W�=��V�4�Q�V�ڗ��`f������Ǘ~�g�7o�<ɧc�]t�c�o~��$u����c�Z[֎���6%����nZS�Ym�M��silu���0 J�ڤbР3)`��W�������Wq=�2K_x�fUs�'k��V��YmE\�A����1z���� }b�4����9�D�	����b��]�E��Ś(���X
p�(eB`��@N
�������%^�+do6W9t+�r�E]Π�������b��kO��Sr�<�?Av=}���Bfݝ㢯vS�L�O�s>���l�$���;T�A7��?O�V�Tl�*�h4�h�d4�W��.��ni[y��dvc2�M��'��]Pe-�o�uf�.�q�!QN�Y��[�/O�Rx���c�!�w1�E;�I� �R����Kkc�-�*Hھ��&���:�N=�{٨���xI��onU�����&�V��qL����76n�M�2�V�u����wT�/�pX���YƯ����eY��b�CX�<�9�q��C�����?=���k�%j��v���s�,�a2j&�Z���H�73�L�SV�p/�fp&V��U7�Э]ߗr�}C1c��*�-�ڹ4�9�&6�2��Xl<�9�Ll��/{�T�9�;G���6���j��q?����2ݨAԴ���@S*��ߥÎɩ�5�7��5N�� M��[[�.պ3���w/��5����:ː�W8�����Օ�<h4- ��`y�N�O[�-�L��p'�-o.ڠ�h�m�v7�ln��ʳ����9޳�?)�ݱ}�^���Gj��2�Ͻ|7;h�	���5�ۅٞu���`E���1�5�F���711�i��5����]kin�(l5`K�{`:�R�N�׵a�G����nMCi���s{2�黯��ۂ��*_1䛸{���ۘϳ:�
���ݜ$���/c����C��짎czcgqrG;o=*��ݽ)+�3�ʄ�	�%$2��ά��э/j"�w^��6FN�+8��������k���~#{�b޿�6Bu�.xTy�b5�h����������;$�P5��U���ɻ�lǶ�y��}j��&���z�����^�uK����F���oS&�y�dZ7���V���i]uf��T�q/��EH5�=.�����L(|I���I�"�6D����2����t`�[�K!&�؄[.^0��tǺ�u,o�46�
�Y'ս�r�=��O��[Yy�^����+������Iݾd�Hod޽�2��&��xh�\��Qt��Xe6�tj�}n�3.o�7�����%�@E�*l�U�����V\�����r ��T&}ld�z�۞:�m	�m���g�xӭ�>��{�Ooz��;�g�ۧݚidN6���zn��� yW��m����ff!Q�+&���ԵU�,�v�S��0:�WJ��{*f�.�ę3p��\�L��,F�s~|���6�|�[��p��<-�r�����M�d&�ky�2:��խF쨝�
̎}.�W@�U�M�1/�_(�\gMv��4��IsZzaڄ���D(I�Caʉ��>G��x�t�[J2��̳�!���P�O8#���+k� �R��ԁ:����꿬T�#�:e��dt*�$�'.Q��߾�M�����;���8Kr{nFVX����F�^W��L�	0�!��h8M�U/�ܘ�&�*��cl]fW�kw����7[~).py߫�1�x5p���3?��	�H���->gs���Cؐ#�K8���J�<��O	~Y=��}�r6����2\���%��P�EK>��!S�<�]��+U	G�SmWwW��/�y��G����z�����L_��T�=i����F��^ò��XEmޘ��k������<p���#��]��-��HA���ʀ`4fﺶn���L���9�a�&�
�U�w?�DW��\Wj����A�u�;�� ���Kxx-�i�SL���b�o���hJ���W��}������U�����U8.≥���"��+�-�E+ Ү5٦���`�3����[�:����<8f_p�(�5�������ݔ-L'�F��h5ަf�f�4-�����N�z�3w��L�t�Ѯ��q��mh��B��ܖ=�M��ͺ{5s:�J4���q�5cw;Y]\Λh��ĳhƕ_q�,m��" W3N,���V;��,?�� NX��������A��h�u��GMB�[���4+�e�I�8�l6���2�M-��2���X�EB�F�6�\�컵���	v3��tك��]U.�\�[0�Q�l���a�7��cfa Yfcٮ�h��.���r2�ZF��P[,�թ�u�3M9gV�0�0����AfvKƗ�B:Lq��pYs��դ���T���@�l������#��]{f���+���͟�uTs	��]5<F�]6�DD�Z�-�T�+�wI��M��WjcmX�팁�mڮ:�hKI���ԯmB55���F��(�%-j�8�*�Sbd6��_�b%~ʉ��h�!������t=�ӆ\KOia�}�r�O�-�b�����+�z|ໆA�>G�)�F�7��mN�喺�����e�a �%���&S.=��](��*f��*5+���ƪ��kxW(�c���B���'��pݬ13q�Sw�4̽7+�d{�`�U�oJ��$e(�]�:)^p�.p����m��Qj�����Ja����_�Cn��}�7�?f�</~T�����
�xv�<����ت���D���o�v�a�}~��o�ǹ�U����=&��������z��!zI:�,�	��0�*�M(C�|�^�&�m��᰷hwt��U{��^�uU�}&0Ol�nײ��%FX�׏��y����=�*}+M��f�FQ�~	�\p�-�*C�Vz�U� \������qQ�UYP/�_�\����T&��H��h�/ ���9�@C����4����)�zm�Ca�K��-��n�·]��&��ǳ6'.k�NTb���'���rOR,;�{��g9l����[�뿣�>b�����Um�ɥ�u��9�]��-�K���`�pS	+)t4Еi䙥q�le;:�:4- SAAl	���w��k�'��{�S6e��,�Nc��炄am�t�bw���-�������,g��(���9e���E��~��X_Dd�&l6�L2KB&�����Kvof�;�G��`C�m+�|FU�%��aB¿uO�}��}����d�7jz���[A��ުz�?���}�YO���b�Y=��<=��^7�|gl��ݰ���$4�4@*%`N�^5�P����b�[���i�M1|5>��Q�?���}B��w��)�9W{  ��o�NL�%�LLRU��zyA�$����ﳓ���ֲ���Q�V�m����XL�@4!�$	���~�U^�D�z}�0�b%�@Lz�.�T�+����(Ue�B"3R���X[.g�/�|�ܝ��'J���X�&D�5�Ȏ��K�#xl_C�8v�Md�4���! ���i8�p����Q�9��P"l�n�/�>s^w��ɥ,�'ʧ����uc�f��'7�7'����!��jNl���Y�*B��=/M(�l�tF�g~��#���<��߷�Ɵej�uf3ql���{9-�,4��k�����x�ecW�S�b�:�%.�K�l%R�`ݖY��׾n��6��o�q�.U��B�l�*�nJH(}���${j>��}��{>�+�7}���L��y\l�]��Շ�Z�����=%��}^P6
E�`6 ���e�ڦ1��۱����v��}�7q?e��.�ͻ�*��t��6�v/3�ŚѬ��m�y�>�ݴ���eq��=83Y�|z�Ƕ�u�;�T�#��$i���V��콌�2q^Q�'�]� ���H"ȇ�̂�A�9f�ֻn�(TׇT���s=�0e<��##5��W# ��%�8�W�p+B����Ą�TЭ�J#}[�Wiٹ}�Y�ו9��ibۄ�4��?��su����䣝2��3F_e5&iTa��]倛��w�*V�J*�� [��G�}1��s�Ogi.���<�;`#�_V�.<]-�yk�����ymq�N�x=��f�$m�ej������R�6��ѝy�&Kn}��Dl�N��^�w��,-Mg��Ң	�U1w��R������u�y�%{/�(�}"
�K �C$��	�*0x�֗ǃ�4��i��lZT�H��y�[�f��7oF�٬���K�_�4�o�9i��<��x�ˊ��'v�֠�Zf��>G����:��������_�~����S;pݲ\E���~�=����_�eF��	!x�x�%毄���#�\Ҫ�V':���Ԝ����"������ꌐ#no�κ�47rgs���왘8:�q�Q3�d8�翳��{�2��
�s�1L��ݪ �1h:�j��9�^�l�c�Z�2�46.KjlZ�q(�o?y�����%���R�qd9����=:Z9"�=��3��Y��񔮵F>~U>5��{�F�f.:���$�S�C�o�R�D����0��AC	�r��m/V�`�I��7~�}�M����(�,�2B�v�'rk��i)'�մр��8��mdb����k�Ѷ{�o�^�fS|�_#_{h��0'qIo���ϧ��¿~'�"�[��:+�������Py<*�kX�=��|;����-�z�{>~�?��B���f�ό�f���I5�i�\�#���\^Ά2�6���m�ݔ�������'Gs�;~�]Uz???g�a���Z�.��[�3��)����/h/��2��ϔ4����ܦq�.����Y���c�xc0�����k�H��W�{fjUrLS���7�צ����3�;�=)!g�o~�~���Yu�(����z�\mi#�$�D0��ʩ>��u[�-�v59٦a��
�ZjM�^��ttl��(�
��v.p�s�cp���������	�����Q���ū�I����1��F�i�7Mq��ЬIM�!i5m)��48�9� �Ah[e2�e��BL7�-�H%��>Cn�uQ>;k����f�@�O�Vܟ�B���Y�ݟG:"�ݹ�!�l&��j�b�jfJ���C�+���3�2[qr�g"��P�|��7��7n��[�/�o������ޅX+"��}����m�E��Gkٮ�]���+T�%M��QE��uyS+�{TSލ����ee�l���n&w�;����{U5��7-I>�/S'/�X\�L�[�[ 8�K� 2�a����A~ָyj����w�{��f���yp�.m����(N�v%��P�Fǃf�s-��}�Z^���W��#��^Y5;�-�!�q�wի���C�W�7�g�@�W8�������<���i{f
h��>���V���̪k�ӡ[�7&��;��n问�CK#ĻZS��վ�v{�ۤ�3f����
�LTbF)�� 'h8 ��%��(!�YbO,�����Sd�tE��=��=�ng�������,���N�h��X%G�]�@�z�k�[���V��h��bVȟ�J��}�Z�-���@����<���Iw9�L��o��B���_�����*��B	%)�@$�����`﭅aH��\�o��YB� ��$�`S�>��z��%�@!���, =dR%@
DT�,�&g�FI	4�I1�(O֬�!��Hߺ�@o(���i	�@0HI� j@����X �O���4��R�A|6z�.�P R�d�I$���*�������a�ݓ�j~�/��V��v'ҩ���Y9Y���l4}Y���H�>j�O���`.��+Ѡ�y>�*�hF���?�Gi����w��@A_�l,d�����?$��2U� /a!�aO�D�/PN���wb��V�!&���	@|�T�pr?�
��J�� ����< ��Ca�3�8���$3}�/Y�	=�� �?N�t͛�uH�¨S=�i���m4�j;:��*Cd �#��~��0�?�~����dX��BҘ*�H�Z�y�7N��EB��C�s6�d�S&��b��9��@��
+&�+,u� �b��w��e���6��m�l��]Ѡ�j��^
����;�G��X��%B
MX θ���'ٵ%4k-[sk+��n���+%@fVk��7�,���g�Lۖ)�nN�O���u^i��0�����xո�H�
ZK��7W���b^	�ܶ�N��);�+kl��l�,�R��4���΄��(*d$0�d@��HRЄ)i	,������ H 2� @@�I��RdŖ�6@m��vT�`E�'��� *�ԅ$������Kp��$�>�n�sJ�[�3�
_�`-2�`S�>~�$ >�]��XA�0Aj��&MɓL�� ����A��^���+�`��
��x��(M�v�N1�����{ã������Iqn'�����D0k�'�~�� ��N�XSQsy�{��,\�e9(+*�����L��c�����)D�AA�K˒�~���h �sa|b0��1[��Fp�5>d	I�VYCs��~����9�`��+e�����w$��ѹ�95�ɠ��B�O�g`!�@AY%B.8��� ��5��y�K��91DU箃7��?�K��@|.6?��a4s�Q����D[��v�Ns��ޅ���c~��Hs����2����g]��=��o�o%4��k��X  �2�q��N���R3�ˌ�=P��&n#����q�o4�ɤ��J���hX/�PV��4�wm%�v��I�BS:H4���f0��s��3n$Op*�$�9�h8
�����X��q$waac���T]��(��pk�T�W<ZI<���T��spR �e2h�+ş�Pa��w$S�	M�ؐ