BZh91AY&SYl� g߀Px����߰����P�[��F�[i��S�Ii�$��)�f���6�j� �5OѠIP        �B)�44�e<�� h�&��@�F&#M0CL�h0	�	�m4SO)�4=5=F@  �JYo���B%$$@�!>��D���RX��BL�[Nj8:( �%f3#����A����m5��Dܲi׮���'��拧�����"����i�xXn4^F@�<zѹ�K��P��*�~șDQHPy���x�pH��<��u�@���+oޕ���  N\T	ht��[ro�9xQߵ�I���Z�����5�U��ϙ.6�ޗ�n5��$܋���T�m���S��Ϛ�䕖h��*���ݠ���J��6��%�p��&��%�5�SY�7X�[ćI�lю�1V\:kqF���`��VK�8l��I �j�2&B�m�N�3I0�N�l���0�����kŒ�n 6���6!9i�L������yȇ����'�%�#CVw��C�Xێk�������O��4��pji���ۧ���~��4�����ߑy|	�Y�JM�G�3M�j�F��c�
	d!8 :���������e�����M2삶M�Z����IY�qT����柨�юܘ�Nyz��]&o	x��/����(���Ѫ��	�p��Ex�A�����x�HA�~zvp��PXz��8ΐ�WǑ�J�CW�y�R�T6�]}"���{t�oD���@H]d�ֻFj٬B\��g���T�RΨ�L�Ø�9���e(�:3�S��{.&~�À��&�x�����Q:婒1�&na#����_�&���"����s���~7P0���f
W@�PK�h�pq.<%�(ce��
򅊅*�S�V}Ld�7ԣ;]V���G!i�\�����e�̳���NS@ �7[i�s:�����3�6��xY͓	 o�K��n�-�G���H+L����*d�xI<�Ԕ�p�����(��H���XP�*���V�*ZA�E6�j�Q �)�9f��k����$	��D������[��兣���2���Z��cI����*�͐!(ѦIFP��`���9�Q�~+�PV�CL
lD�2����ʇ���ۘ��T^A��N�I��#�EAYL�!,a%ӄ��-��BRb@��F22�Q��q��[e
1.˖4� �TĲ(p�J����b�U�X��e^r�k�i��W���e�eR������d�4��a���H�
m�P@